(0 + 0) => x"37", (0 + 1) => x"41", (0 + 2) => x"00", (0 + 3) => x"00", (0 + 4) => x"6f", (0 + 5) => x"00", (0 + 6) => x"60", (0 + 7) => x"2f", (0 + 8) => x"79", (0 + 9) => x"71", (0 + 10) => x"1c", (0 + 11) => x"08", (0 + 12) => x"11", (0 + 13) => x"6e", (0 + 14) => x"22", (0 + 15) => x"d6", (0 + 16) => x"26", (0 + 17) => x"d4", (0 + 18) => x"4a", (0 + 19) => x"d2", (0 + 20) => x"4e", (0 + 21) => x"d0", (0 + 22) => x"33", (0 + 23) => x"86", (0 + 24) => x"c7", (0 + 25) => x"01", (0 + 26) => x"52", (0 + 27) => x"ce", (0 + 28) => x"56", (0 + 29) => x"cc", (0 + 30) => x"5a", (0 + 31) => x"ca", (0 + 32) => x"91", (0 + 33) => x"67", (0 + 34) => x"23", (0 + 35) => x"80", (0 + 36) => x"07", (0 + 37) => x"00", (0 + 38) => x"97", (0 + 39) => x"08", (0 + 40) => x"00", (0 + 41) => x"00", (0 + 42) => x"93", (0 + 43) => x"88", (0 + 44) => x"68", (0 + 45) => x"65", (0 + 46) => x"17", (0 + 47) => x"04", (0 + 48) => x"00", (0 + 49) => x"00", (0 + 50) => x"13", (0 + 51) => x"04", (0 + 52) => x"64", (0 + 53) => x"64", (0 + 54) => x"01", (0 + 55) => x"43", (0 + 56) => x"81", (0 + 57) => x"4e", (0 + 58) => x"29", (0 + 59) => x"4f", (0 + 60) => x"05", (0 + 61) => x"47", (0 + 62) => x"cd", (0 + 63) => x"45", (0 + 64) => x"d5", (0 + 65) => x"46", (0 + 66) => x"39", (0 + 67) => x"16", (0 + 68) => x"ad", (0 + 69) => x"43", (0 + 70) => x"31", (0 + 71) => x"68", (0 + 72) => x"93", (0 + 73) => x"02", (0 + 74) => x"f0", (0 + 75) => x"03", (0 + 76) => x"c1", (0 + 77) => x"6f", (0 + 78) => x"fd", (0 + 79) => x"59", (0 + 80) => x"21", (0 + 81) => x"49", (0 + 82) => x"85", (0 + 83) => x"44", (0 + 84) => x"97", (0 + 85) => x"47", (0 + 86) => x"00", (0 + 87) => x"00", (0 + 88) => x"23", (0 + 89) => x"88", (0 + 90) => x"e7", (0 + 91) => x"62", (0 + 92) => x"97", (0 + 93) => x"47", (0 + 94) => x"00", (0 + 95) => x"00", (0 + 96) => x"23", (0 + 97) => x"8c", (0 + 98) => x"e7", (0 + 99) => x"60", (0 + 100) => x"03", (0 + 101) => x"2a", (0 + 102) => x"05", (0 + 103) => x"00", (0 + 104) => x"97", (0 + 105) => x"07", (0 + 106) => x"00", (0 + 107) => x"00", (0 + 108) => x"93", (0 + 109) => x"87", (0 + 110) => x"c7", (0 + 111) => x"60", (0 + 112) => x"72", (0 + 113) => x"9a", (0 + 114) => x"23", (0 + 115) => x"00", (0 + 116) => x"ea", (0 + 117) => x"00", (0 + 118) => x"85", (0 + 119) => x"07", (0 + 120) => x"03", (0 + 121) => x"ca", (0 + 122) => x"07", (0 + 123) => x"00", (0 + 124) => x"e3", (0 + 125) => x"1d", (0 + 126) => x"0a", (0 + 127) => x"fe", (0 + 128) => x"03", (0 + 129) => x"2a", (0 + 130) => x"05", (0 + 131) => x"00", (0 + 132) => x"81", (0 + 133) => x"8f", (0 + 134) => x"83", (0 + 135) => x"4a", (0 + 136) => x"0a", (0 + 137) => x"00", (0 + 138) => x"52", (0 + 139) => x"8b", (0 + 140) => x"63", (0 + 141) => x"81", (0 + 142) => x"0a", (0 + 143) => x"14", (0 + 144) => x"05", (0 + 145) => x"0a", (0 + 146) => x"83", (0 + 147) => x"4a", (0 + 148) => x"0a", (0 + 149) => x"00", (0 + 150) => x"e3", (0 + 151) => x"9d", (0 + 152) => x"0a", (0 + 153) => x"fe", (0 + 154) => x"33", (0 + 155) => x"0a", (0 + 156) => x"6a", (0 + 157) => x"41", (0 + 158) => x"8d", (0 + 159) => x"07", (0 + 160) => x"d2", (0 + 161) => x"97", (0 + 162) => x"13", (0 + 163) => x"8a", (0 + 164) => x"17", (0 + 165) => x"00", (0 + 166) => x"63", (0 + 167) => x"e9", (0 + 168) => x"f5", (0 + 169) => x"00", (0 + 170) => x"97", (0 + 171) => x"47", (0 + 172) => x"00", (0 + 173) => x"00", (0 + 174) => x"23", (0 + 175) => x"8d", (0 + 176) => x"e7", (0 + 177) => x"5e", (0 + 178) => x"05", (0 + 179) => x"0a", (0 + 180) => x"e3", (0 + 181) => x"1b", (0 + 182) => x"da", (0 + 183) => x"fe", (0 + 184) => x"97", (0 + 185) => x"47", (0 + 186) => x"00", (0 + 187) => x"00", (0 + 188) => x"23", (0 + 189) => x"88", (0 + 190) => x"e7", (0 + 191) => x"5c", (0 + 192) => x"97", (0 + 193) => x"47", (0 + 194) => x"00", (0 + 195) => x"00", (0 + 196) => x"23", (0 + 197) => x"82", (0 + 198) => x"e7", (0 + 199) => x"5c", (0 + 200) => x"97", (0 + 201) => x"47", (0 + 202) => x"00", (0 + 203) => x"00", (0 + 204) => x"23", (0 + 205) => x"8a", (0 + 206) => x"e7", (0 + 207) => x"5a", (0 + 208) => x"93", (0 + 209) => x"07", (0 + 210) => x"e1", (0 + 211) => x"00", (0 + 212) => x"f2", (0 + 213) => x"97", (0 + 214) => x"23", (0 + 215) => x"80", (0 + 216) => x"e7", (0 + 217) => x"00", (0 + 218) => x"f9", (0 + 219) => x"17", (0 + 220) => x"e3", (0 + 221) => x"1d", (0 + 222) => x"f6", (0 + 223) => x"fe", (0 + 224) => x"97", (0 + 225) => x"07", (0 + 226) => x"00", (0 + 227) => x"00", (0 + 228) => x"93", (0 + 229) => x"87", (0 + 230) => x"c7", (0 + 231) => x"59", (0 + 232) => x"85", (0 + 233) => x"07", (0 + 234) => x"03", (0 + 235) => x"ca", (0 + 236) => x"07", (0 + 237) => x"00", (0 + 238) => x"e3", (0 + 239) => x"1d", (0 + 240) => x"0a", (0 + 241) => x"fe", (0 + 242) => x"b3", (0 + 243) => x"87", (0 + 244) => x"17", (0 + 245) => x"41", (0 + 246) => x"13", (0 + 247) => x"8a", (0 + 248) => x"b7", (0 + 249) => x"00", (0 + 250) => x"b1", (0 + 251) => x"07", (0 + 252) => x"63", (0 + 253) => x"e9", (0 + 254) => x"45", (0 + 255) => x"01", (0 + 256) => x"17", (0 + 257) => x"4a", (0 + 258) => x"00", (0 + 259) => x"00", (0 + 260) => x"23", (0 + 261) => x"02", (0 + 262) => x"ea", (0 + 263) => x"5a", (0 + 264) => x"85", (0 + 265) => x"07", (0 + 266) => x"e3", (0 + 267) => x"9b", (0 + 268) => x"d7", (0 + 269) => x"fe", (0 + 270) => x"97", (0 + 271) => x"07", (0 + 272) => x"00", (0 + 273) => x"00", (0 + 274) => x"93", (0 + 275) => x"87", (0 + 276) => x"e7", (0 + 277) => x"56", (0 + 278) => x"85", (0 + 279) => x"07", (0 + 280) => x"03", (0 + 281) => x"ca", (0 + 282) => x"07", (0 + 283) => x"00", (0 + 284) => x"e3", (0 + 285) => x"1d", (0 + 286) => x"0a", (0 + 287) => x"fe", (0 + 288) => x"b3", (0 + 289) => x"87", (0 + 290) => x"17", (0 + 291) => x"41", (0 + 292) => x"b3", (0 + 293) => x"07", (0 + 294) => x"ff", (0 + 295) => x"40", (0 + 296) => x"13", (0 + 297) => x"8a", (0 + 298) => x"17", (0 + 299) => x"00", (0 + 300) => x"63", (0 + 301) => x"e9", (0 + 302) => x"f5", (0 + 303) => x"00", (0 + 304) => x"97", (0 + 305) => x"47", (0 + 306) => x"00", (0 + 307) => x"00", (0 + 308) => x"23", (0 + 309) => x"8a", (0 + 310) => x"e7", (0 + 311) => x"56", (0 + 312) => x"05", (0 + 313) => x"0a", (0 + 314) => x"e3", (0 + 315) => x"1b", (0 + 316) => x"da", (0 + 317) => x"fe", (0 + 318) => x"97", (0 + 319) => x"47", (0 + 320) => x"00", (0 + 321) => x"00", (0 + 322) => x"23", (0 + 323) => x"81", (0 + 324) => x"e7", (0 + 325) => x"56", (0 + 326) => x"97", (0 + 327) => x"07", (0 + 328) => x"00", (0 + 329) => x"00", (0 + 330) => x"93", (0 + 331) => x"87", (0 + 332) => x"67", (0 + 333) => x"53", (0 + 334) => x"85", (0 + 335) => x"07", (0 + 336) => x"03", (0 + 337) => x"ca", (0 + 338) => x"07", (0 + 339) => x"00", (0 + 340) => x"e3", (0 + 341) => x"1d", (0 + 342) => x"0a", (0 + 343) => x"fe", (0 + 344) => x"33", (0 + 345) => x"8a", (0 + 346) => x"63", (0 + 347) => x"40", (0 + 348) => x"b3", (0 + 349) => x"87", (0 + 350) => x"17", (0 + 351) => x"41", (0 + 352) => x"d2", (0 + 353) => x"97", (0 + 354) => x"13", (0 + 355) => x"8a", (0 + 356) => x"17", (0 + 357) => x"00", (0 + 358) => x"63", (0 + 359) => x"e9", (0 + 360) => x"f5", (0 + 361) => x"00", (0 + 362) => x"97", (0 + 363) => x"47", (0 + 364) => x"00", (0 + 365) => x"00", (0 + 366) => x"23", (0 + 367) => x"8d", (0 + 368) => x"e7", (0 + 369) => x"52", (0 + 370) => x"05", (0 + 371) => x"0a", (0 + 372) => x"e3", (0 + 373) => x"1b", (0 + 374) => x"da", (0 + 375) => x"fe", (0 + 376) => x"23", (0 + 377) => x"11", (0 + 378) => x"58", (0 + 379) => x"00", (0 + 380) => x"23", (0 + 381) => x"02", (0 + 382) => x"08", (0 + 383) => x"00", (0 + 384) => x"83", (0 + 385) => x"57", (0 + 386) => x"08", (0 + 387) => x"00", (0 + 388) => x"23", (0 + 389) => x"80", (0 + 390) => x"0f", (0 + 391) => x"00", (0 + 392) => x"c2", (0 + 393) => x"07", (0 + 394) => x"c1", (0 + 395) => x"83", (0 + 396) => x"13", (0 + 397) => x"fa", (0 + 398) => x"17", (0 + 399) => x"00", (0 + 400) => x"63", (0 + 401) => x"09", (0 + 402) => x"0a", (0 + 403) => x"00", (0 + 404) => x"93", (0 + 405) => x"17", (0 + 406) => x"43", (0 + 407) => x"00", (0 + 408) => x"b3", (0 + 409) => x"97", (0 + 410) => x"f4", (0 + 411) => x"00", (0 + 412) => x"b3", (0 + 413) => x"8e", (0 + 414) => x"fe", (0 + 415) => x"40", (0 + 416) => x"55", (0 + 417) => x"bd", (0 + 418) => x"13", (0 + 419) => x"fa", (0 + 420) => x"27", (0 + 421) => x"00", (0 + 422) => x"63", (0 + 423) => x"08", (0 + 424) => x"0a", (0 + 425) => x"00", (0 + 426) => x"93", (0 + 427) => x"17", (0 + 428) => x"43", (0 + 429) => x"00", (0 + 430) => x"b3", (0 + 431) => x"97", (0 + 432) => x"f4", (0 + 433) => x"00", (0 + 434) => x"be", (0 + 435) => x"9e", (0 + 436) => x"45", (0 + 437) => x"b5", (0 + 438) => x"13", (0 + 439) => x"ff", (0 + 440) => x"07", (0 + 441) => x"01", (0 + 442) => x"63", (0 + 443) => x"0c", (0 + 444) => x"0f", (0 + 445) => x"00", (0 + 446) => x"05", (0 + 447) => x"03", (0 + 448) => x"13", (0 + 449) => x"0f", (0 + 450) => x"a3", (0 + 451) => x"00", (0 + 452) => x"e3", (0 + 453) => x"18", (0 + 454) => x"23", (0 + 455) => x"e9", (0 + 456) => x"01", (0 + 457) => x"43", (0 + 458) => x"29", (0 + 459) => x"4f", (0 + 460) => x"61", (0 + 461) => x"b5", (0 + 462) => x"01", (0 + 463) => x"4a", (0 + 464) => x"f9", (0 + 465) => x"b5", (0 + 466) => x"13", (0 + 467) => x"ff", (0 + 468) => x"07", (0 + 469) => x"02", (0 + 470) => x"63", (0 + 471) => x"0a", (0 + 472) => x"0f", (0 + 473) => x"00", (0 + 474) => x"7d", (0 + 475) => x"13", (0 + 476) => x"13", (0 + 477) => x"0f", (0 + 478) => x"a3", (0 + 479) => x"00", (0 + 480) => x"e3", (0 + 481) => x"1a", (0 + 482) => x"33", (0 + 483) => x"e7", (0 + 484) => x"1d", (0 + 485) => x"43", (0 + 486) => x"45", (0 + 487) => x"4f", (0 + 488) => x"b5", (0 + 489) => x"b5", (0 + 490) => x"91", (0 + 491) => x"8b", (0 + 492) => x"81", (0 + 493) => x"c7", (0 + 494) => x"5c", (0 + 495) => x"41", (0 + 496) => x"23", (0 + 497) => x"a0", (0 + 498) => x"d7", (0 + 499) => x"01", (0 + 500) => x"32", (0 + 501) => x"54", (0 + 502) => x"a2", (0 + 503) => x"54", (0 + 504) => x"12", (0 + 505) => x"59", (0 + 506) => x"82", (0 + 507) => x"59", (0 + 508) => x"72", (0 + 509) => x"4a", (0 + 510) => x"e2", (0 + 511) => x"4a", (0 + 512) => x"52", (0 + 513) => x"4b", (0 + 514) => x"45", (0 + 515) => x"61", (0 + 516) => x"82", (0 + 517) => x"80", (0 + 518) => x"91", (0 + 519) => x"65", (0 + 520) => x"23", (0 + 521) => x"80", (0 + 522) => x"05", (0 + 523) => x"00", (0 + 524) => x"85", (0 + 525) => x"46", (0 + 526) => x"97", (0 + 527) => x"47", (0 + 528) => x"00", (0 + 529) => x"00", (0 + 530) => x"23", (0 + 531) => x"8b", (0 + 532) => x"d7", (0 + 533) => x"46", (0 + 534) => x"97", (0 + 535) => x"47", (0 + 536) => x"00", (0 + 537) => x"00", (0 + 538) => x"23", (0 + 539) => x"89", (0 + 540) => x"d7", (0 + 541) => x"48", (0 + 542) => x"18", (0 + 543) => x"41", (0 + 544) => x"17", (0 + 545) => x"06", (0 + 546) => x"00", (0 + 547) => x"00", (0 + 548) => x"13", (0 + 549) => x"06", (0 + 550) => x"86", (0 + 551) => x"48", (0 + 552) => x"41", (0 + 553) => x"11", (0 + 554) => x"2e", (0 + 555) => x"97", (0 + 556) => x"b2", (0 + 557) => x"87", (0 + 558) => x"23", (0 + 559) => x"00", (0 + 560) => x"d7", (0 + 561) => x"00", (0 + 562) => x"85", (0 + 563) => x"07", (0 + 564) => x"03", (0 + 565) => x"c7", (0 + 566) => x"07", (0 + 567) => x"00", (0 + 568) => x"6d", (0 + 569) => x"ff", (0 + 570) => x"18", (0 + 571) => x"41", (0 + 572) => x"91", (0 + 573) => x"8f", (0 + 574) => x"83", (0 + 575) => x"46", (0 + 576) => x"07", (0 + 577) => x"00", (0 + 578) => x"3a", (0 + 579) => x"86", (0 + 580) => x"cd", (0 + 581) => x"ca", (0 + 582) => x"05", (0 + 583) => x"07", (0 + 584) => x"83", (0 + 585) => x"46", (0 + 586) => x"07", (0 + 587) => x"00", (0 + 588) => x"ed", (0 + 589) => x"fe", (0 + 590) => x"11", (0 + 591) => x"8f", (0 + 592) => x"8d", (0 + 593) => x"07", (0 + 594) => x"ba", (0 + 595) => x"97", (0 + 596) => x"cd", (0 + 597) => x"46", (0 + 598) => x"13", (0 + 599) => x"87", (0 + 600) => x"17", (0 + 601) => x"00", (0 + 602) => x"63", (0 + 603) => x"eb", (0 + 604) => x"f6", (0 + 605) => x"00", (0 + 606) => x"85", (0 + 607) => x"46", (0 + 608) => x"d5", (0 + 609) => x"47", (0 + 610) => x"17", (0 + 611) => x"46", (0 + 612) => x"00", (0 + 613) => x"00", (0 + 614) => x"23", (0 + 615) => x"01", (0 + 616) => x"d6", (0 + 617) => x"44", (0 + 618) => x"05", (0 + 619) => x"07", (0 + 620) => x"e3", (0 + 621) => x"1b", (0 + 622) => x"f7", (0 + 623) => x"fe", (0 + 624) => x"85", (0 + 625) => x"46", (0 + 626) => x"17", (0 + 627) => x"47", (0 + 628) => x"00", (0 + 629) => x"00", (0 + 630) => x"23", (0 + 631) => x"0b", (0 + 632) => x"d7", (0 + 633) => x"40", (0 + 634) => x"17", (0 + 635) => x"47", (0 + 636) => x"00", (0 + 637) => x"00", (0 + 638) => x"23", (0 + 639) => x"05", (0 + 640) => x"d7", (0 + 641) => x"40", (0 + 642) => x"91", (0 + 643) => x"67", (0 + 644) => x"18", (0 + 645) => x"08", (0 + 646) => x"3e", (0 + 647) => x"97", (0 + 648) => x"17", (0 + 649) => x"46", (0 + 650) => x"00", (0 + 651) => x"00", (0 + 652) => x"23", (0 + 653) => x"0a", (0 + 654) => x"d6", (0 + 655) => x"3e", (0 + 656) => x"93", (0 + 657) => x"06", (0 + 658) => x"e1", (0 + 659) => x"00", (0 + 660) => x"b6", (0 + 661) => x"97", (0 + 662) => x"39", (0 + 663) => x"17", (0 + 664) => x"85", (0 + 665) => x"46", (0 + 666) => x"23", (0 + 667) => x"80", (0 + 668) => x"d7", (0 + 669) => x"00", (0 + 670) => x"f9", (0 + 671) => x"17", (0 + 672) => x"e3", (0 + 673) => x"1d", (0 + 674) => x"f7", (0 + 675) => x"fe", (0 + 676) => x"97", (0 + 677) => x"06", (0 + 678) => x"00", (0 + 679) => x"00", (0 + 680) => x"93", (0 + 681) => x"86", (0 + 682) => x"86", (0 + 683) => x"3d", (0 + 684) => x"b6", (0 + 685) => x"87", (0 + 686) => x"85", (0 + 687) => x"07", (0 + 688) => x"03", (0 + 689) => x"c7", (0 + 690) => x"07", (0 + 691) => x"00", (0 + 692) => x"6d", (0 + 693) => x"ff", (0 + 694) => x"95", (0 + 695) => x"8f", (0 + 696) => x"93", (0 + 697) => x"86", (0 + 698) => x"b7", (0 + 699) => x"00", (0 + 700) => x"4d", (0 + 701) => x"47", (0 + 702) => x"b1", (0 + 703) => x"07", (0 + 704) => x"63", (0 + 705) => x"6b", (0 + 706) => x"d7", (0 + 707) => x"00", (0 + 708) => x"85", (0 + 709) => x"46", (0 + 710) => x"55", (0 + 711) => x"47", (0 + 712) => x"17", (0 + 713) => x"46", (0 + 714) => x"00", (0 + 715) => x"00", (0 + 716) => x"23", (0 + 717) => x"0e", (0 + 718) => x"d6", (0 + 719) => x"3c", (0 + 720) => x"85", (0 + 721) => x"07", (0 + 722) => x"e3", (0 + 723) => x"9b", (0 + 724) => x"e7", (0 + 725) => x"fe", (0 + 726) => x"85", (0 + 727) => x"47", (0 + 728) => x"17", (0 + 729) => x"47", (0 + 730) => x"00", (0 + 731) => x"00", (0 + 732) => x"23", (0 + 733) => x"08", (0 + 734) => x"f7", (0 + 735) => x"3a", (0 + 736) => x"21", (0 + 737) => x"47", (0 + 738) => x"b1", (0 + 739) => x"67", (0 + 740) => x"23", (0 + 741) => x"91", (0 + 742) => x"e7", (0 + 743) => x"00", (0 + 744) => x"23", (0 + 745) => x"82", (0 + 746) => x"07", (0 + 747) => x"00", (0 + 748) => x"c1", (0 + 749) => x"67", (0 + 750) => x"23", (0 + 751) => x"80", (0 + 752) => x"07", (0 + 753) => x"00", (0 + 754) => x"41", (0 + 755) => x"01", (0 + 756) => x"82", (0 + 757) => x"80", (0 + 758) => x"01", (0 + 759) => x"47", (0 + 760) => x"a1", (0 + 761) => x"bf", (0 + 762) => x"17", (0 + 763) => x"27", (0 + 764) => x"00", (0 + 765) => x"00", (0 + 766) => x"23", (0 + 767) => x"23", (0 + 768) => x"07", (0 + 769) => x"d0", (0 + 770) => x"37", (0 + 771) => x"57", (0 + 772) => x"34", (0 + 773) => x"12", (0 + 774) => x"35", (0 + 775) => x"71", (0 + 776) => x"97", (0 + 777) => x"07", (0 + 778) => x"00", (0 + 779) => x"00", (0 + 780) => x"93", (0 + 781) => x"87", (0 + 782) => x"87", (0 + 783) => x"39", (0 + 784) => x"13", (0 + 785) => x"07", (0 + 786) => x"87", (0 + 787) => x"67", (0 + 788) => x"97", (0 + 789) => x"26", (0 + 790) => x"00", (0 + 791) => x"00", (0 + 792) => x"23", (0 + 793) => x"a8", (0 + 794) => x"e6", (0 + 795) => x"ce", (0 + 796) => x"3e", (0 + 797) => x"c6", (0 + 798) => x"3e", (0 + 799) => x"c8", (0 + 800) => x"3e", (0 + 801) => x"ca", (0 + 802) => x"97", (0 + 803) => x"07", (0 + 804) => x"00", (0 + 805) => x"00", (0 + 806) => x"93", (0 + 807) => x"87", (0 + 808) => x"27", (0 + 809) => x"38", (0 + 810) => x"06", (0 + 811) => x"cf", (0 + 812) => x"22", (0 + 813) => x"cd", (0 + 814) => x"26", (0 + 815) => x"cb", (0 + 816) => x"4a", (0 + 817) => x"c9", (0 + 818) => x"4e", (0 + 819) => x"c7", (0 + 820) => x"52", (0 + 821) => x"c5", (0 + 822) => x"56", (0 + 823) => x"c3", (0 + 824) => x"5a", (0 + 825) => x"c1", (0 + 826) => x"de", (0 + 827) => x"de", (0 + 828) => x"e2", (0 + 829) => x"dc", (0 + 830) => x"e6", (0 + 831) => x"da", (0 + 832) => x"3e", (0 + 833) => x"cc", (0 + 834) => x"01", (0 + 835) => x"47", (0 + 836) => x"13", (0 + 837) => x"06", (0 + 838) => x"80", (0 + 839) => x"05", (0 + 840) => x"93", (0 + 841) => x"06", (0 + 842) => x"00", (0 + 843) => x"02", (0 + 844) => x"d1", (0 + 845) => x"48", (0 + 846) => x"9c", (0 + 847) => x"18", (0 + 848) => x"ba", (0 + 849) => x"97", (0 + 850) => x"23", (0 + 851) => x"86", (0 + 852) => x"c7", (0 + 853) => x"fa", (0 + 854) => x"a3", (0 + 855) => x"80", (0 + 856) => x"c7", (0 + 857) => x"fc", (0 + 858) => x"93", (0 + 859) => x"05", (0 + 860) => x"17", (0 + 861) => x"00", (0 + 862) => x"23", (0 + 863) => x"8b", (0 + 864) => x"c7", (0 + 865) => x"fc", (0 + 866) => x"13", (0 + 867) => x"88", (0 + 868) => x"15", (0 + 869) => x"00", (0 + 870) => x"13", (0 + 871) => x"85", (0 + 872) => x"25", (0 + 873) => x"00", (0 + 874) => x"a3", (0 + 875) => x"85", (0 + 876) => x"c7", (0 + 877) => x"fe", (0 + 878) => x"0d", (0 + 879) => x"8b", (0 + 880) => x"13", (0 + 881) => x"f3", (0 + 882) => x"35", (0 + 883) => x"00", (0 + 884) => x"13", (0 + 885) => x"78", (0 + 886) => x"38", (0 + 887) => x"00", (0 + 888) => x"0d", (0 + 889) => x"89", (0 + 890) => x"19", (0 + 891) => x"e3", (0 + 892) => x"23", (0 + 893) => x"86", (0 + 894) => x"d7", (0 + 895) => x"fa", (0 + 896) => x"63", (0 + 897) => x"14", (0 + 898) => x"03", (0 + 899) => x"00", (0 + 900) => x"a3", (0 + 901) => x"80", (0 + 902) => x"d7", (0 + 903) => x"fc", (0 + 904) => x"63", (0 + 905) => x"14", (0 + 906) => x"08", (0 + 907) => x"00", (0 + 908) => x"23", (0 + 909) => x"8b", (0 + 910) => x"d7", (0 + 911) => x"fc", (0 + 912) => x"19", (0 + 913) => x"e1", (0 + 914) => x"a3", (0 + 915) => x"85", (0 + 916) => x"d7", (0 + 917) => x"fe", (0 + 918) => x"2e", (0 + 919) => x"87", (0 + 920) => x"e3", (0 + 921) => x"9b", (0 + 922) => x"15", (0 + 923) => x"fb", (0 + 924) => x"23", (0 + 925) => x"08", (0 + 926) => x"01", (0 + 927) => x"02", (0 + 928) => x"a3", (0 + 929) => x"02", (0 + 930) => x"01", (0 + 931) => x"04", (0 + 932) => x"23", (0 + 933) => x"0d", (0 + 934) => x"01", (0 + 935) => x"04", (0 + 936) => x"a3", (0 + 937) => x"07", (0 + 938) => x"01", (0 + 939) => x"06", (0 + 940) => x"91", (0 + 941) => x"67", (0 + 942) => x"23", (0 + 943) => x"80", (0 + 944) => x"07", (0 + 945) => x"00", (0 + 946) => x"85", (0 + 947) => x"67", (0 + 948) => x"31", (0 + 949) => x"67", (0 + 950) => x"93", (0 + 951) => x"87", (0 + 952) => x"07", (0 + 953) => x"80", (0 + 954) => x"23", (0 + 955) => x"11", (0 + 956) => x"f7", (0 + 957) => x"00", (0 + 958) => x"13", (0 + 959) => x"07", (0 + 960) => x"40", (0 + 961) => x"1f", (0 + 962) => x"a1", (0 + 963) => x"67", (0 + 964) => x"23", (0 + 965) => x"90", (0 + 966) => x"e7", (0 + 967) => x"00", (0 + 968) => x"21", (0 + 969) => x"4e", (0 + 970) => x"05", (0 + 971) => x"46", (0 + 972) => x"89", (0 + 973) => x"48", (0 + 974) => x"05", (0 + 975) => x"48", (0 + 976) => x"0d", (0 + 977) => x"45", (0 + 978) => x"81", (0 + 979) => x"46", (0 + 980) => x"a1", (0 + 981) => x"6f", (0 + 982) => x"91", (0 + 983) => x"65", (0 + 984) => x"05", (0 + 985) => x"47", (0 + 986) => x"7d", (0 + 987) => x"5f", (0 + 988) => x"b1", (0 + 989) => x"6e", (0 + 990) => x"13", (0 + 991) => x"93", (0 + 992) => x"26", (0 + 993) => x"00", (0 + 994) => x"b3", (0 + 995) => x"07", (0 + 996) => x"d3", (0 + 997) => x"00", (0 + 998) => x"80", (0 + 999) => x"18", (0 + 1000) => x"23", (0 + 1001) => x"81", (0 + 1002) => x"0f", (0 + 1003) => x"00", (0 + 1004) => x"22", (0 + 1005) => x"93", (0 + 1006) => x"8a", (0 + 1007) => x"07", (0 + 1008) => x"b6", (0 + 1009) => x"97", (0 + 1010) => x"83", (0 + 1011) => x"22", (0 + 1012) => x"c3", (0 + 1013) => x"f9", (0 + 1014) => x"60", (0 + 1015) => x"08", (0 + 1016) => x"a2", (0 + 1017) => x"97", (0 + 1018) => x"13", (0 + 1019) => x"13", (0 + 1020) => x"25", (0 + 1021) => x"00", (0 + 1022) => x"80", (0 + 1023) => x"18", (0 + 1024) => x"ae", (0 + 1025) => x"97", (0 + 1026) => x"23", (0 + 1027) => x"80", (0 + 1028) => x"e7", (0 + 1029) => x"00", (0 + 1030) => x"22", (0 + 1031) => x"93", (0 + 1032) => x"93", (0 + 1033) => x"17", (0 + 1034) => x"28", (0 + 1035) => x"00", (0 + 1036) => x"ae", (0 + 1037) => x"92", (0 + 1038) => x"23", (0 + 1039) => x"80", (0 + 1040) => x"e2", (0 + 1041) => x"00", (0 + 1042) => x"a2", (0 + 1043) => x"97", (0 + 1044) => x"83", (0 + 1045) => x"23", (0 + 1046) => x"c3", (0 + 1047) => x"f9", (0 + 1048) => x"17", (0 + 1049) => x"44", (0 + 1050) => x"00", (0 + 1051) => x"00", (0 + 1052) => x"23", (0 + 1053) => x"06", (0 + 1054) => x"e4", (0 + 1055) => x"26", (0 + 1056) => x"83", (0 + 1057) => x"a2", (0 + 1058) => x"c7", (0 + 1059) => x"f9", (0 + 1060) => x"80", (0 + 1061) => x"18", (0 + 1062) => x"97", (0 + 1063) => x"47", (0 + 1064) => x"00", (0 + 1065) => x"00", (0 + 1066) => x"23", (0 + 1067) => x"8b", (0 + 1068) => x"e7", (0 + 1069) => x"28", (0 + 1070) => x"13", (0 + 1071) => x"93", (0 + 1072) => x"28", (0 + 1073) => x"00", (0 + 1074) => x"22", (0 + 1075) => x"93", (0 + 1076) => x"ae", (0 + 1077) => x"93", (0 + 1078) => x"17", (0 + 1079) => x"44", (0 + 1080) => x"00", (0 + 1081) => x"00", (0 + 1082) => x"23", (0 + 1083) => x"01", (0 + 1084) => x"e4", (0 + 1085) => x"26", (0 + 1086) => x"23", (0 + 1087) => x"80", (0 + 1088) => x"e3", (0 + 1089) => x"00", (0 + 1090) => x"93", (0 + 1091) => x"17", (0 + 1092) => x"26", (0 + 1093) => x"00", (0 + 1094) => x"ae", (0 + 1095) => x"92", (0 + 1096) => x"23", (0 + 1097) => x"80", (0 + 1098) => x"e2", (0 + 1099) => x"00", (0 + 1100) => x"b2", (0 + 1101) => x"97", (0 + 1102) => x"03", (0 + 1103) => x"23", (0 + 1104) => x"c3", (0 + 1105) => x"f9", (0 + 1106) => x"17", (0 + 1107) => x"44", (0 + 1108) => x"00", (0 + 1109) => x"00", (0 + 1110) => x"23", (0 + 1111) => x"0b", (0 + 1112) => x"e4", (0 + 1113) => x"26", (0 + 1114) => x"8a", (0 + 1115) => x"07", (0 + 1116) => x"b2", (0 + 1117) => x"97", (0 + 1118) => x"60", (0 + 1119) => x"08", (0 + 1120) => x"2e", (0 + 1121) => x"93", (0 + 1122) => x"a2", (0 + 1123) => x"97", (0 + 1124) => x"93", (0 + 1125) => x"83", (0 + 1126) => x"d6", (0 + 1127) => x"ff", (0 + 1128) => x"23", (0 + 1129) => x"00", (0 + 1130) => x"e3", (0 + 1131) => x"00", (0 + 1132) => x"ae", (0 + 1133) => x"97", (0 + 1134) => x"05", (0 + 1135) => x"05", (0 + 1136) => x"05", (0 + 1137) => x"08", (0 + 1138) => x"85", (0 + 1139) => x"08", (0 + 1140) => x"b3", (0 + 1141) => x"33", (0 + 1142) => x"70", (0 + 1143) => x"00", (0 + 1144) => x"23", (0 + 1145) => x"80", (0 + 1146) => x"e7", (0 + 1147) => x"00", (0 + 1148) => x"93", (0 + 1149) => x"02", (0 + 1150) => x"c5", (0 + 1151) => x"ff", (0 + 1152) => x"13", (0 + 1153) => x"03", (0 + 1154) => x"c8", (0 + 1155) => x"ff", (0 + 1156) => x"93", (0 + 1157) => x"87", (0 + 1158) => x"c8", (0 + 1159) => x"ff", (0 + 1160) => x"85", (0 + 1161) => x"06", (0 + 1162) => x"b3", (0 + 1163) => x"03", (0 + 1164) => x"70", (0 + 1165) => x"40", (0 + 1166) => x"b3", (0 + 1167) => x"32", (0 + 1168) => x"50", (0 + 1169) => x"00", (0 + 1170) => x"33", (0 + 1171) => x"33", (0 + 1172) => x"60", (0 + 1173) => x"00", (0 + 1174) => x"b3", (0 + 1175) => x"37", (0 + 1176) => x"f0", (0 + 1177) => x"00", (0 + 1178) => x"7d", (0 + 1179) => x"16", (0 + 1180) => x"7d", (0 + 1181) => x"1e", (0 + 1182) => x"b3", (0 + 1183) => x"02", (0 + 1184) => x"50", (0 + 1185) => x"40", (0 + 1186) => x"33", (0 + 1187) => x"03", (0 + 1188) => x"60", (0 + 1189) => x"40", (0 + 1190) => x"b3", (0 + 1191) => x"07", (0 + 1192) => x"f0", (0 + 1193) => x"40", (0 + 1194) => x"b3", (0 + 1195) => x"f6", (0 + 1196) => x"76", (0 + 1197) => x"00", (0 + 1198) => x"63", (0 + 1199) => x"13", (0 + 1200) => x"e6", (0 + 1201) => x"01", (0 + 1202) => x"0d", (0 + 1203) => x"46", (0 + 1204) => x"23", (0 + 1205) => x"82", (0 + 1206) => x"0e", (0 + 1207) => x"00", (0 + 1208) => x"33", (0 + 1209) => x"75", (0 + 1210) => x"55", (0 + 1211) => x"00", (0 + 1212) => x"33", (0 + 1213) => x"78", (0 + 1214) => x"68", (0 + 1215) => x"00", (0 + 1216) => x"b3", (0 + 1217) => x"f8", (0 + 1218) => x"f8", (0 + 1219) => x"00", (0 + 1220) => x"e3", (0 + 1221) => x"1d", (0 + 1222) => x"0e", (0 + 1223) => x"f0", (0 + 1224) => x"97", (0 + 1225) => x"0c", (0 + 1226) => x"00", (0 + 1227) => x"00", (0 + 1228) => x"93", (0 + 1229) => x"8c", (0 + 1230) => x"8c", (0 + 1231) => x"1e", (0 + 1232) => x"13", (0 + 1233) => x"0c", (0 + 1234) => x"40", (0 + 1235) => x"60", (0 + 1236) => x"91", (0 + 1237) => x"6b", (0 + 1238) => x"05", (0 + 1239) => x"44", (0 + 1240) => x"cd", (0 + 1241) => x"44", (0 + 1242) => x"91", (0 + 1243) => x"49", (0 + 1244) => x"23", (0 + 1245) => x"80", (0 + 1246) => x"0b", (0 + 1247) => x"00", (0 + 1248) => x"09", (0 + 1249) => x"4b", (0 + 1250) => x"81", (0 + 1251) => x"4a", (0 + 1252) => x"01", (0 + 1253) => x"4a", (0 + 1254) => x"55", (0 + 1255) => x"49", (0 + 1256) => x"97", (0 + 1257) => x"47", (0 + 1258) => x"00", (0 + 1259) => x"00", (0 + 1260) => x"23", (0 + 1261) => x"8e", (0 + 1262) => x"87", (0 + 1263) => x"18", (0 + 1264) => x"97", (0 + 1265) => x"47", (0 + 1266) => x"00", (0 + 1267) => x"00", (0 + 1268) => x"23", (0 + 1269) => x"80", (0 + 1270) => x"87", (0 + 1271) => x"1c", (0 + 1272) => x"97", (0 + 1273) => x"07", (0 + 1274) => x"00", (0 + 1275) => x"00", (0 + 1276) => x"93", (0 + 1277) => x"87", (0 + 1278) => x"87", (0 + 1279) => x"1b", (0 + 1280) => x"85", (0 + 1281) => x"07", (0 + 1282) => x"03", (0 + 1283) => x"c7", (0 + 1284) => x"07", (0 + 1285) => x"00", (0 + 1286) => x"6d", (0 + 1287) => x"ff", (0 + 1288) => x"b3", (0 + 1289) => x"87", (0 + 1290) => x"97", (0 + 1291) => x"41", (0 + 1292) => x"13", (0 + 1293) => x"87", (0 + 1294) => x"37", (0 + 1295) => x"00", (0 + 1296) => x"91", (0 + 1297) => x"07", (0 + 1298) => x"63", (0 + 1299) => x"e9", (0 + 1300) => x"e4", (0 + 1301) => x"00", (0 + 1302) => x"17", (0 + 1303) => x"47", (0 + 1304) => x"00", (0 + 1305) => x"00", (0 + 1306) => x"23", (0 + 1307) => x"07", (0 + 1308) => x"87", (0 + 1309) => x"18", (0 + 1310) => x"85", (0 + 1311) => x"07", (0 + 1312) => x"e3", (0 + 1313) => x"9b", (0 + 1314) => x"27", (0 + 1315) => x"ff", (0 + 1316) => x"63", (0 + 1317) => x"44", (0 + 1318) => x"5b", (0 + 1319) => x"03", (0 + 1320) => x"13", (0 + 1321) => x"96", (0 + 1322) => x"1a", (0 + 1323) => x"00", (0 + 1324) => x"56", (0 + 1325) => x"96", (0 + 1326) => x"0a", (0 + 1327) => x"06", (0 + 1328) => x"62", (0 + 1329) => x"96", (0 + 1330) => x"13", (0 + 1331) => x"05", (0 + 1332) => x"1b", (0 + 1333) => x"00", (0 + 1334) => x"56", (0 + 1335) => x"87", (0 + 1336) => x"63", (0 + 1337) => x"d3", (0 + 1338) => x"e9", (0 + 1339) => x"04", (0 + 1340) => x"97", (0 + 1341) => x"47", (0 + 1342) => x"00", (0 + 1343) => x"00", (0 + 1344) => x"23", (0 + 1345) => x"86", (0 + 1346) => x"87", (0 + 1347) => x"14", (0 + 1348) => x"05", (0 + 1349) => x"07", (0 + 1350) => x"31", (0 + 1351) => x"06", (0 + 1352) => x"e3", (0 + 1353) => x"18", (0 + 1354) => x"a7", (0 + 1355) => x"fe", (0 + 1356) => x"b1", (0 + 1357) => x"67", (0 + 1358) => x"3d", (0 + 1359) => x"47", (0 + 1360) => x"23", (0 + 1361) => x"91", (0 + 1362) => x"e7", (0 + 1363) => x"00", (0 + 1364) => x"23", (0 + 1365) => x"82", (0 + 1366) => x"07", (0 + 1367) => x"00", (0 + 1368) => x"83", (0 + 1369) => x"d7", (0 + 1370) => x"07", (0 + 1371) => x"00", (0 + 1372) => x"41", (0 + 1373) => x"67", (0 + 1374) => x"23", (0 + 1375) => x"00", (0 + 1376) => x"07", (0 + 1377) => x"00", (0 + 1378) => x"c2", (0 + 1379) => x"07", (0 + 1380) => x"c1", (0 + 1381) => x"83", (0 + 1382) => x"13", (0 + 1383) => x"f7", (0 + 1384) => x"17", (0 + 1385) => x"00", (0 + 1386) => x"31", (0 + 1387) => x"cf", (0 + 1388) => x"8d", (0 + 1389) => x"47", (0 + 1390) => x"e3", (0 + 1391) => x"cd", (0 + 1392) => x"47", (0 + 1393) => x"f7", (0 + 1394) => x"05", (0 + 1395) => x"0a", (0 + 1396) => x"e3", (0 + 1397) => x"5a", (0 + 1398) => x"4b", (0 + 1399) => x"f7", (0 + 1400) => x"85", (0 + 1401) => x"0a", (0 + 1402) => x"05", (0 + 1403) => x"0b", (0 + 1404) => x"b5", (0 + 1405) => x"b7", (0 + 1406) => x"63", (0 + 1407) => x"0d", (0 + 1408) => x"47", (0 + 1409) => x"07", (0 + 1410) => x"97", (0 + 1411) => x"47", (0 + 1412) => x"00", (0 + 1413) => x"00", (0 + 1414) => x"23", (0 + 1415) => x"81", (0 + 1416) => x"87", (0 + 1417) => x"10", (0 + 1418) => x"1c", (0 + 1419) => x"42", (0 + 1420) => x"de", (0 + 1421) => x"97", (0 + 1422) => x"23", (0 + 1423) => x"80", (0 + 1424) => x"87", (0 + 1425) => x"00", (0 + 1426) => x"0c", (0 + 1427) => x"42", (0 + 1428) => x"83", (0 + 1429) => x"c7", (0 + 1430) => x"05", (0 + 1431) => x"00", (0 + 1432) => x"b1", (0 + 1433) => x"c3", (0 + 1434) => x"ae", (0 + 1435) => x"87", (0 + 1436) => x"85", (0 + 1437) => x"07", (0 + 1438) => x"83", (0 + 1439) => x"c6", (0 + 1440) => x"07", (0 + 1441) => x"00", (0 + 1442) => x"ed", (0 + 1443) => x"fe", (0 + 1444) => x"8d", (0 + 1445) => x"8f", (0 + 1446) => x"93", (0 + 1447) => x"86", (0 + 1448) => x"37", (0 + 1449) => x"00", (0 + 1450) => x"91", (0 + 1451) => x"07", (0 + 1452) => x"63", (0 + 1453) => x"f4", (0 + 1454) => x"d4", (0 + 1455) => x"00", (0 + 1456) => x"51", (0 + 1457) => x"bf", (0 + 1458) => x"b6", (0 + 1459) => x"87", (0 + 1460) => x"97", (0 + 1461) => x"46", (0 + 1462) => x"00", (0 + 1463) => x"00", (0 + 1464) => x"23", (0 + 1465) => x"88", (0 + 1466) => x"86", (0 + 1467) => x"0e", (0 + 1468) => x"93", (0 + 1469) => x"86", (0 + 1470) => x"17", (0 + 1471) => x"00", (0 + 1472) => x"e3", (0 + 1473) => x"f9", (0 + 1474) => x"f4", (0 + 1475) => x"fe", (0 + 1476) => x"41", (0 + 1477) => x"b7", (0 + 1478) => x"13", (0 + 1479) => x"f7", (0 + 1480) => x"27", (0 + 1481) => x"00", (0 + 1482) => x"19", (0 + 1483) => x"cb", (0 + 1484) => x"e3", (0 + 1485) => x"0e", (0 + 1486) => x"0a", (0 + 1487) => x"f0", (0 + 1488) => x"7d", (0 + 1489) => x"1a", (0 + 1490) => x"e3", (0 + 1491) => x"5b", (0 + 1492) => x"5a", (0 + 1493) => x"f1", (0 + 1494) => x"fd", (0 + 1495) => x"1a", (0 + 1496) => x"7d", (0 + 1497) => x"1b", (0 + 1498) => x"39", (0 + 1499) => x"b7", (0 + 1500) => x"91", (0 + 1501) => x"47", (0 + 1502) => x"d9", (0 + 1503) => x"bf", (0 + 1504) => x"91", (0 + 1505) => x"8b", (0 + 1506) => x"e3", (0 + 1507) => x"8d", (0 + 1508) => x"07", (0 + 1509) => x"ee", (0 + 1510) => x"93", (0 + 1511) => x"17", (0 + 1512) => x"1a", (0 + 1513) => x"00", (0 + 1514) => x"d2", (0 + 1515) => x"97", (0 + 1516) => x"8a", (0 + 1517) => x"07", (0 + 1518) => x"e2", (0 + 1519) => x"97", (0 + 1520) => x"d8", (0 + 1521) => x"43", (0 + 1522) => x"88", (0 + 1523) => x"47", (0 + 1524) => x"02", (0 + 1525) => x"97", (0 + 1526) => x"cd", (0 + 1527) => x"bd", (0 + 1528) => x"97", (0 + 1529) => x"47", (0 + 1530) => x"00", (0 + 1531) => x"00", (0 + 1532) => x"23", (0 + 1533) => x"82", (0 + 1534) => x"87", (0 + 1535) => x"0e", (0 + 1536) => x"69", (0 + 1537) => x"b7", (0 + 1538) => x"00", (0 + 1539) => x"00", (0 + 1540) => x"e0", (0 + 1541) => x"06", (0 + 1542) => x"00", (0 + 1543) => x"00", (0 + 1544) => x"06", (0 + 1545) => x"02", (0 + 1546) => x"00", (0 + 1547) => x"00", (0 + 1548) => x"5c", (0 + 1549) => x"06", (0 + 1550) => x"00", (0 + 1551) => x"00", (0 + 1552) => x"f4", (0 + 1553) => x"06", (0 + 1554) => x"00", (0 + 1555) => x"00", (0 + 1556) => x"06", (0 + 1557) => x"02", (0 + 1558) => x"00", (0 + 1559) => x"00", (0 + 1560) => x"64", (0 + 1561) => x"06", (0 + 1562) => x"00", (0 + 1563) => x"00", (0 + 1564) => x"08", (0 + 1565) => x"07", (0 + 1566) => x"00", (0 + 1567) => x"00", (0 + 1568) => x"08", (0 + 1569) => x"00", (0 + 1570) => x"00", (0 + 1571) => x"00", (0 + 1572) => x"64", (0 + 1573) => x"06", (0 + 1574) => x"00", (0 + 1575) => x"00", (0 + 1576) => x"1c", (0 + 1577) => x"07", (0 + 1578) => x"00", (0 + 1579) => x"00", (0 + 1580) => x"06", (0 + 1581) => x"02", (0 + 1582) => x"00", (0 + 1583) => x"00", (0 + 1584) => x"6c", (0 + 1585) => x"06", (0 + 1586) => x"00", (0 + 1587) => x"00", (0 + 1588) => x"30", (0 + 1589) => x"07", (0 + 1590) => x"00", (0 + 1591) => x"00", (0 + 1592) => x"08", (0 + 1593) => x"00", (0 + 1594) => x"00", (0 + 1595) => x"00", (0 + 1596) => x"6c", (0 + 1597) => x"06", (0 + 1598) => x"00", (0 + 1599) => x"00", (0 + 1600) => x"30", (0 + 1601) => x"31", (0 + 1602) => x"32", (0 + 1603) => x"33", (0 + 1604) => x"34", (0 + 1605) => x"35", (0 + 1606) => x"36", (0 + 1607) => x"37", (0 + 1608) => x"38", (0 + 1609) => x"39", (0 + 1610) => x"41", (0 + 1611) => x"42", (0 + 1612) => x"43", (0 + 1613) => x"44", (0 + 1614) => x"45", (0 + 1615) => x"46", (0 + 1616) => x"b0", (0 + 1617) => x"06", (0 + 1618) => x"00", (0 + 1619) => x"00", (0 + 1620) => x"04", (0 + 1621) => x"06", (0 + 1622) => x"00", (0 + 1623) => x"00", (0 + 1624) => x"05", (0 + 1625) => x"00", (0 + 1626) => x"00", (0 + 1627) => x"00", (0 + 1628) => x"e8", (0 + 1629) => x"06", (0 + 1630) => x"00", (0 + 1631) => x"00", (0 + 1632) => x"44", (0 + 1633) => x"07", (0 + 1634) => x"00", (0 + 1635) => x"00", (0 + 1636) => x"10", (0 + 1637) => x"07", (0 + 1638) => x"00", (0 + 1639) => x"00", (0 + 1640) => x"00", (0 + 1641) => x"20", (0 + 1642) => x"00", (0 + 1643) => x"00", (0 + 1644) => x"38", (0 + 1645) => x"07", (0 + 1646) => x"00", (0 + 1647) => x"00", (0 + 1648) => x"04", (0 + 1649) => x"20", (0 + 1650) => x"00", (0 + 1651) => x"00", (0 + 1652) => x"53", (0 + 1653) => x"45", (0 + 1654) => x"54", (0 + 1655) => x"20", (0 + 1656) => x"20", (0 + 1657) => x"3a", (0 + 1658) => x"20", (0 + 1659) => x"00", (0 + 1660) => x"56", (0 + 1661) => x"41", (0 + 1662) => x"4c", (0 + 1663) => x"55", (0 + 1664) => x"45", (0 + 1665) => x"3a", (0 + 1666) => x"20", (0 + 1667) => x"00", (0 + 1668) => x"20", (0 + 1669) => x"20", (0 + 1670) => x"20", (0 + 1671) => x"00", (0 + 1672) => x"20", (0 + 1673) => x"20", (0 + 1674) => x"20", (0 + 1675) => x"20", (0 + 1676) => x"20", (0 + 1677) => x"20", (0 + 1678) => x"20", (0 + 1679) => x"20", (0 + 1680) => x"20", (0 + 1681) => x"20", (0 + 1682) => x"20", (0 + 1683) => x"20", (0 + 1684) => x"20", (0 + 1685) => x"20", (0 + 1686) => x"20", (0 + 1687) => x"20", (0 + 1688) => x"20", (0 + 1689) => x"20", (0 + 1690) => x"20", (0 + 1691) => x"20", (0 + 1692) => x"00", (0 + 1693) => x"00", (0 + 1694) => x"00", (0 + 1695) => x"00", (0 + 1696) => x"58", (0 + 1697) => x"00", (0 + 1698) => x"00", (0 + 1699) => x"00", (0 + 1700) => x"20", (0 + 1701) => x"00", (0 + 1702) => x"00", (0 + 1703) => x"00", (0 + 1704) => x"4e", (0 + 1705) => x"41", (0 + 1706) => x"4d", (0 + 1707) => x"45", (0 + 1708) => x"20", (0 + 1709) => x"3a", (0 + 1710) => x"20", (0 + 1711) => x"00", (0 + 1712) => x"4d", (0 + 1713) => x"41", (0 + 1714) => x"49", (0 + 1715) => x"4e", (0 + 1716) => x"20", (0 + 1717) => x"4d", (0 + 1718) => x"45", (0 + 1719) => x"4e", (0 + 1720) => x"55", (0 + 1721) => x"00", (0 + 1722) => x"00", (0 + 1723) => x"00", (0 + 1724) => x"53", (0 + 1725) => x"54", (0 + 1726) => x"41", (0 + 1727) => x"52", (0 + 1728) => x"54", (0 + 1729) => x"49", (0 + 1730) => x"4e", (0 + 1731) => x"47", (0 + 1732) => x"20", (0 + 1733) => x"55", (0 + 1734) => x"50", (0 + 1735) => x"00", (0 + 1736) => x"20", (0 + 1737) => x"20", (0 + 1738) => x"20", (0 + 1739) => x"20", (0 + 1740) => x"20", (0 + 1741) => x"20", (0 + 1742) => x"20", (0 + 1743) => x"20", (0 + 1744) => x"20", (0 + 1745) => x"20", (0 + 1746) => x"20", (0 + 1747) => x"20", (0 + 1748) => x"20", (0 + 1749) => x"20", (0 + 1750) => x"20", (0 + 1751) => x"20", (0 + 1752) => x"20", (0 + 1753) => x"20", (0 + 1754) => x"00", (0 + 1755) => x"00", (0 + 1756) => x"20", (0 + 1757) => x"58", (0 + 1758) => x"20", (0 + 1759) => x"00", (0 + 1760) => x"31", (0 + 1761) => x"2e", (0 + 1762) => x"20", (0 + 1763) => x"73", (0 + 1764) => x"68", (0 + 1765) => x"6f", (0 + 1766) => x"77", (0 + 1767) => x"20", (0 + 1768) => x"6d", (0 + 1769) => x"79", (0 + 1770) => x"5f", (0 + 1771) => x"76", (0 + 1772) => x"61", (0 + 1773) => x"6c", (0 + 1774) => x"5f", (0 + 1775) => x"72", (0 + 1776) => x"6f", (0 + 1777) => x"6d", (0 + 1778) => x"00", (0 + 1779) => x"00", (0 + 1780) => x"32", (0 + 1781) => x"2e", (0 + 1782) => x"20", (0 + 1783) => x"73", (0 + 1784) => x"68", (0 + 1785) => x"6f", (0 + 1786) => x"77", (0 + 1787) => x"20", (0 + 1788) => x"6d", (0 + 1789) => x"79", (0 + 1790) => x"5f", (0 + 1791) => x"76", (0 + 1792) => x"61", (0 + 1793) => x"6c", (0 + 1794) => x"5f", (0 + 1795) => x"72", (0 + 1796) => x"61", (0 + 1797) => x"6d", (0 + 1798) => x"31", (0 + 1799) => x"00", (0 + 1800) => x"33", (0 + 1801) => x"2e", (0 + 1802) => x"20", (0 + 1803) => x"73", (0 + 1804) => x"65", (0 + 1805) => x"74", (0 + 1806) => x"20", (0 + 1807) => x"20", (0 + 1808) => x"6d", (0 + 1809) => x"79", (0 + 1810) => x"5f", (0 + 1811) => x"76", (0 + 1812) => x"61", (0 + 1813) => x"6c", (0 + 1814) => x"5f", (0 + 1815) => x"72", (0 + 1816) => x"61", (0 + 1817) => x"6d", (0 + 1818) => x"31", (0 + 1819) => x"00", (0 + 1820) => x"34", (0 + 1821) => x"2e", (0 + 1822) => x"20", (0 + 1823) => x"73", (0 + 1824) => x"68", (0 + 1825) => x"6f", (0 + 1826) => x"77", (0 + 1827) => x"20", (0 + 1828) => x"6d", (0 + 1829) => x"79", (0 + 1830) => x"5f", (0 + 1831) => x"76", (0 + 1832) => x"61", (0 + 1833) => x"6c", (0 + 1834) => x"5f", (0 + 1835) => x"72", (0 + 1836) => x"61", (0 + 1837) => x"6d", (0 + 1838) => x"32", (0 + 1839) => x"00", (0 + 1840) => x"35", (0 + 1841) => x"2e", (0 + 1842) => x"20", (0 + 1843) => x"73", (0 + 1844) => x"65", (0 + 1845) => x"74", (0 + 1846) => x"20", (0 + 1847) => x"20", (0 + 1848) => x"6d", (0 + 1849) => x"79", (0 + 1850) => x"5f", (0 + 1851) => x"76", (0 + 1852) => x"61", (0 + 1853) => x"6c", (0 + 1854) => x"5f", (0 + 1855) => x"72", (0 + 1856) => x"61", (0 + 1857) => x"6d", (0 + 1858) => x"32", (0 + 1859) => x"00", (0 + 1860) => x"ef", (0 + 1861) => x"be", (0 + 1862) => x"ad", (0 + 1863) => x"de", (0 + 1864) => x"00", (0 + 1865) => x"00", (0 + 1866) => x"00", (0 + 1867) => x"00", (0 + 1868) => x"00", (0 + 1869) => x"00", (0 + 1870) => x"00", (0 + 1871) => x"00", (0 + 1872) => x"00", (0 + 1873) => x"00", (0 + 1874) => x"00", (0 + 1875) => x"00", (0 + 1876) => x"00", (0 + 1877) => x"00", (0 + 1878) => x"00", (0 + 1879) => x"00", (0 + 1880) => x"00", (0 + 1881) => x"00", (0 + 1882) => x"00", (0 + 1883) => x"00", (0 + 1884) => x"00", (0 + 1885) => x"00", (0 + 1886) => x"00", (0 + 1887) => x"00", (0 + 1888) => x"00", (0 + 1889) => x"00", (0 + 1890) => x"00", (0 + 1891) => x"00", (0 + 1892) => x"00", (0 + 1893) => x"00", (0 + 1894) => x"00", (0 + 1895) => x"00", (0 + 1896) => x"00", (0 + 1897) => x"00", (0 + 1898) => x"00", (0 + 1899) => x"00", (0 + 1900) => x"00", (0 + 1901) => x"00", (0 + 1902) => x"00", (0 + 1903) => x"00", (0 + 1904) => x"00", (0 + 1905) => x"00", (0 + 1906) => x"00", (0 + 1907) => x"00", (0 + 1908) => x"00", (0 + 1909) => x"00", (0 + 1910) => x"00", (0 + 1911) => x"00", (0 + 1912) => x"00", (0 + 1913) => x"00", (0 + 1914) => x"00", (0 + 1915) => x"00", (0 + 1916) => x"00", (0 + 1917) => x"00", (0 + 1918) => x"00", (0 + 1919) => x"00", (0 + 1920) => x"00", (0 + 1921) => x"00", (0 + 1922) => x"00", (0 + 1923) => x"00", (0 + 1924) => x"00", (0 + 1925) => x"00", (0 + 1926) => x"00", (0 + 1927) => x"00", (0 + 1928) => x"00", (0 + 1929) => x"00", (0 + 1930) => x"00", (0 + 1931) => x"00", (0 + 1932) => x"00", (0 + 1933) => x"00", (0 + 1934) => x"00", (0 + 1935) => x"00", (0 + 1936) => x"00", (0 + 1937) => x"00", (0 + 1938) => x"00", (0 + 1939) => x"00", (0 + 1940) => x"00", (0 + 1941) => x"00", (0 + 1942) => x"00", (0 + 1943) => x"00", (0 + 1944) => x"00", (0 + 1945) => x"00", (0 + 1946) => x"00", (0 + 1947) => x"00", (0 + 1948) => x"00", (0 + 1949) => x"00", (0 + 1950) => x"00", (0 + 1951) => x"00", (0 + 1952) => x"00", (0 + 1953) => x"00", (0 + 1954) => x"00", (0 + 1955) => x"00", (0 + 1956) => x"00", (0 + 1957) => x"00", (0 + 1958) => x"00", (0 + 1959) => x"00", (0 + 1960) => x"00", (0 + 1961) => x"00", (0 + 1962) => x"00", (0 + 1963) => x"00", (0 + 1964) => x"00", (0 + 1965) => x"00", (0 + 1966) => x"00", (0 + 1967) => x"00", (0 + 1968) => x"00", (0 + 1969) => x"00", (0 + 1970) => x"00", (0 + 1971) => x"00", (0 + 1972) => x"00", (0 + 1973) => x"00", (0 + 1974) => x"00", (0 + 1975) => x"00", (0 + 1976) => x"00", (0 + 1977) => x"00", (0 + 1978) => x"00", (0 + 1979) => x"00", (0 + 1980) => x"00", (0 + 1981) => x"00", (0 + 1982) => x"00", (0 + 1983) => x"00", (0 + 1984) => x"00", (0 + 1985) => x"00", (0 + 1986) => x"00", (0 + 1987) => x"00", (0 + 1988) => x"00", (0 + 1989) => x"00", (0 + 1990) => x"00", (0 + 1991) => x"00", (0 + 1992) => x"00", (0 + 1993) => x"00", (0 + 1994) => x"00", (0 + 1995) => x"00", (0 + 1996) => x"00", (0 + 1997) => x"00", (0 + 1998) => x"00", (0 + 1999) => x"00", (0 + 2000) => x"00", (0 + 2001) => x"00", (0 + 2002) => x"00", (0 + 2003) => x"00", (0 + 2004) => x"00", (0 + 2005) => x"00", (0 + 2006) => x"00", (0 + 2007) => x"00", (0 + 2008) => x"00", (0 + 2009) => x"00", (0 + 2010) => x"00", (0 + 2011) => x"00", (0 + 2012) => x"00", (0 + 2013) => x"00", (0 + 2014) => x"00", (0 + 2015) => x"00", (0 + 2016) => x"00", (0 + 2017) => x"00", (0 + 2018) => x"00", (0 + 2019) => x"00", (0 + 2020) => x"00", (0 + 2021) => x"00", (0 + 2022) => x"00", (0 + 2023) => x"00", (0 + 2024) => x"00", (0 + 2025) => x"00", (0 + 2026) => x"00", (0 + 2027) => x"00", (0 + 2028) => x"00", (0 + 2029) => x"00", (0 + 2030) => x"00", (0 + 2031) => x"00", (0 + 2032) => x"00", (0 + 2033) => x"00", (0 + 2034) => x"00", (0 + 2035) => x"00", (0 + 2036) => x"00", (0 + 2037) => x"00", (0 + 2038) => x"00", (0 + 2039) => x"00", (0 + 2040) => x"00", (0 + 2041) => x"00", (0 + 2042) => x"00", (0 + 2043) => x"00", (0 + 2044) => x"00", (0 + 2045) => x"00", (0 + 2046) => x"00", (0 + 2047) => x"00", (0 + 2048) => x"00", (0 + 2049) => x"00", (0 + 2050) => x"00", (0 + 2051) => x"00", (0 + 2052) => x"00", (0 + 2053) => x"00", (0 + 2054) => x"00", (0 + 2055) => x"00", (0 + 2056) => x"00", (0 + 2057) => x"00", (0 + 2058) => x"00", (0 + 2059) => x"00", (0 + 2060) => x"00", (0 + 2061) => x"00", (0 + 2062) => x"00", (0 + 2063) => x"00", (0 + 2064) => x"00", (0 + 2065) => x"00", (0 + 2066) => x"00", (0 + 2067) => x"00", (0 + 2068) => x"00", (0 + 2069) => x"00", (0 + 2070) => x"00", (0 + 2071) => x"00", (0 + 2072) => x"00", (0 + 2073) => x"00", (0 + 2074) => x"00", (0 + 2075) => x"00", (0 + 2076) => x"00", (0 + 2077) => x"00", (0 + 2078) => x"00", (0 + 2079) => x"00", (0 + 2080) => x"00", (0 + 2081) => x"00", (0 + 2082) => x"00", (0 + 2083) => x"00", (0 + 2084) => x"00", (0 + 2085) => x"00", (0 + 2086) => x"00", (0 + 2087) => x"00", (0 + 2088) => x"00", (0 + 2089) => x"00", (0 + 2090) => x"00", (0 + 2091) => x"00", (0 + 2092) => x"00", (0 + 2093) => x"00", (0 + 2094) => x"00", (0 + 2095) => x"00", (0 + 2096) => x"00", (0 + 2097) => x"00", (0 + 2098) => x"00", (0 + 2099) => x"00", (0 + 2100) => x"00", (0 + 2101) => x"00", (0 + 2102) => x"00", (0 + 2103) => x"00", (0 + 2104) => x"00", (0 + 2105) => x"00", (0 + 2106) => x"00", (0 + 2107) => x"00", (0 + 2108) => x"00", (0 + 2109) => x"00", (0 + 2110) => x"00", (0 + 2111) => x"00", (0 + 2112) => x"00", (0 + 2113) => x"00", (0 + 2114) => x"00", (0 + 2115) => x"00", (0 + 2116) => x"00", (0 + 2117) => x"00", (0 + 2118) => x"00", (0 + 2119) => x"00", (0 + 2120) => x"00", (0 + 2121) => x"00", (0 + 2122) => x"00", (0 + 2123) => x"00", (0 + 2124) => x"00", (0 + 2125) => x"00", (0 + 2126) => x"00", (0 + 2127) => x"00", (0 + 2128) => x"00", (0 + 2129) => x"00", (0 + 2130) => x"00", (0 + 2131) => x"00", (0 + 2132) => x"00", (0 + 2133) => x"00", (0 + 2134) => x"00", (0 + 2135) => x"00", (0 + 2136) => x"00", (0 + 2137) => x"00", (0 + 2138) => x"00", (0 + 2139) => x"00", (0 + 2140) => x"00", (0 + 2141) => x"00", (0 + 2142) => x"00", (0 + 2143) => x"00", (0 + 2144) => x"00", (0 + 2145) => x"00", (0 + 2146) => x"00", (0 + 2147) => x"00", (0 + 2148) => x"00", (0 + 2149) => x"00", (0 + 2150) => x"00", (0 + 2151) => x"00", (0 + 2152) => x"00", (0 + 2153) => x"00", (0 + 2154) => x"00", (0 + 2155) => x"00", (0 + 2156) => x"00", (0 + 2157) => x"00", (0 + 2158) => x"00", (0 + 2159) => x"00", (0 + 2160) => x"00", (0 + 2161) => x"00", (0 + 2162) => x"00", (0 + 2163) => x"00", (0 + 2164) => x"00", (0 + 2165) => x"00", (0 + 2166) => x"00", (0 + 2167) => x"00", (0 + 2168) => x"00", (0 + 2169) => x"00", (0 + 2170) => x"00", (0 + 2171) => x"00", (0 + 2172) => x"00", (0 + 2173) => x"00", (0 + 2174) => x"00", (0 + 2175) => x"00", (0 + 2176) => x"00", (0 + 2177) => x"00", (0 + 2178) => x"00", (0 + 2179) => x"00", (0 + 2180) => x"00", (0 + 2181) => x"00", (0 + 2182) => x"00", (0 + 2183) => x"00", (0 + 2184) => x"00", (0 + 2185) => x"00", (0 + 2186) => x"00", (0 + 2187) => x"00", (0 + 2188) => x"00", (0 + 2189) => x"00", (0 + 2190) => x"00", (0 + 2191) => x"00", (0 + 2192) => x"00", (0 + 2193) => x"00", (0 + 2194) => x"00", (0 + 2195) => x"00", (0 + 2196) => x"00", (0 + 2197) => x"00", (0 + 2198) => x"00", (0 + 2199) => x"00", (0 + 2200) => x"00", (0 + 2201) => x"00", (0 + 2202) => x"00", (0 + 2203) => x"00", (0 + 2204) => x"00", (0 + 2205) => x"00", (0 + 2206) => x"00", (0 + 2207) => x"00", (0 + 2208) => x"00", (0 + 2209) => x"00", (0 + 2210) => x"00", (0 + 2211) => x"00", (0 + 2212) => x"00", (0 + 2213) => x"00", (0 + 2214) => x"00", (0 + 2215) => x"00", (0 + 2216) => x"00", (0 + 2217) => x"00", (0 + 2218) => x"00", (0 + 2219) => x"00", (0 + 2220) => x"00", (0 + 2221) => x"00", (0 + 2222) => x"00", (0 + 2223) => x"00", (0 + 2224) => x"00", (0 + 2225) => x"00", (0 + 2226) => x"00", (0 + 2227) => x"00", (0 + 2228) => x"00", (0 + 2229) => x"00", (0 + 2230) => x"00", (0 + 2231) => x"00", (0 + 2232) => x"00", (0 + 2233) => x"00", (0 + 2234) => x"00", (0 + 2235) => x"00", (0 + 2236) => x"00", (0 + 2237) => x"00", (0 + 2238) => x"00", (0 + 2239) => x"00", (0 + 2240) => x"00", (0 + 2241) => x"00", (0 + 2242) => x"00", (0 + 2243) => x"00", (0 + 2244) => x"00", (0 + 2245) => x"00", (0 + 2246) => x"00", (0 + 2247) => x"00", (0 + 2248) => x"00", (0 + 2249) => x"00", (0 + 2250) => x"00", (0 + 2251) => x"00", (0 + 2252) => x"00", (0 + 2253) => x"00", (0 + 2254) => x"00", (0 + 2255) => x"00", (0 + 2256) => x"00", (0 + 2257) => x"00", (0 + 2258) => x"00", (0 + 2259) => x"00", (0 + 2260) => x"00", (0 + 2261) => x"00", (0 + 2262) => x"00", (0 + 2263) => x"00", (0 + 2264) => x"00", (0 + 2265) => x"00", (0 + 2266) => x"00", (0 + 2267) => x"00", (0 + 2268) => x"00", (0 + 2269) => x"00", (0 + 2270) => x"00", (0 + 2271) => x"00", (0 + 2272) => x"00", (0 + 2273) => x"00", (0 + 2274) => x"00", (0 + 2275) => x"00", (0 + 2276) => x"00", (0 + 2277) => x"00", (0 + 2278) => x"00", (0 + 2279) => x"00", (0 + 2280) => x"00", (0 + 2281) => x"00", (0 + 2282) => x"00", (0 + 2283) => x"00", (0 + 2284) => x"00", (0 + 2285) => x"00", (0 + 2286) => x"00", (0 + 2287) => x"00", (0 + 2288) => x"00", (0 + 2289) => x"00", (0 + 2290) => x"00", (0 + 2291) => x"00", (0 + 2292) => x"00", (0 + 2293) => x"00", (0 + 2294) => x"00", (0 + 2295) => x"00", (0 + 2296) => x"00", (0 + 2297) => x"00", (0 + 2298) => x"00", (0 + 2299) => x"00", (0 + 2300) => x"00", (0 + 2301) => x"00", (0 + 2302) => x"00", (0 + 2303) => x"00", (0 + 2304) => x"00", (0 + 2305) => x"00", (0 + 2306) => x"00", (0 + 2307) => x"00", (0 + 2308) => x"00", (0 + 2309) => x"00", (0 + 2310) => x"00", (0 + 2311) => x"00", (0 + 2312) => x"00", (0 + 2313) => x"00", (0 + 2314) => x"00", (0 + 2315) => x"00", (0 + 2316) => x"00", (0 + 2317) => x"00", (0 + 2318) => x"00", (0 + 2319) => x"00", (0 + 2320) => x"00", (0 + 2321) => x"00", (0 + 2322) => x"00", (0 + 2323) => x"00", (0 + 2324) => x"00", (0 + 2325) => x"00", (0 + 2326) => x"00", (0 + 2327) => x"00", (0 + 2328) => x"00", (0 + 2329) => x"00", (0 + 2330) => x"00", (0 + 2331) => x"00", (0 + 2332) => x"00", (0 + 2333) => x"00", (0 + 2334) => x"00", (0 + 2335) => x"00", (0 + 2336) => x"00", (0 + 2337) => x"00", (0 + 2338) => x"00", (0 + 2339) => x"00", (0 + 2340) => x"00", (0 + 2341) => x"00", (0 + 2342) => x"00", (0 + 2343) => x"00", (0 + 2344) => x"00", (0 + 2345) => x"00", (0 + 2346) => x"00", (0 + 2347) => x"00", (0 + 2348) => x"00", (0 + 2349) => x"00", (0 + 2350) => x"00", (0 + 2351) => x"00", (0 + 2352) => x"00", (0 + 2353) => x"00", (0 + 2354) => x"00", (0 + 2355) => x"00", (0 + 2356) => x"00", (0 + 2357) => x"00", (0 + 2358) => x"00", (0 + 2359) => x"00", (0 + 2360) => x"00", (0 + 2361) => x"00", (0 + 2362) => x"00", (0 + 2363) => x"00", (0 + 2364) => x"00", (0 + 2365) => x"00", (0 + 2366) => x"00", (0 + 2367) => x"00", (0 + 2368) => x"00", (0 + 2369) => x"00", (0 + 2370) => x"00", (0 + 2371) => x"00", (0 + 2372) => x"00", (0 + 2373) => x"00", (0 + 2374) => x"00", (0 + 2375) => x"00", (0 + 2376) => x"00", (0 + 2377) => x"00", (0 + 2378) => x"00", (0 + 2379) => x"00", (0 + 2380) => x"00", (0 + 2381) => x"00", (0 + 2382) => x"00", (0 + 2383) => x"00", (0 + 2384) => x"00", (0 + 2385) => x"00", (0 + 2386) => x"00", (0 + 2387) => x"00", (0 + 2388) => x"00", (0 + 2389) => x"00", (0 + 2390) => x"00", (0 + 2391) => x"00", (0 + 2392) => x"00", (0 + 2393) => x"00", (0 + 2394) => x"00", (0 + 2395) => x"00", (0 + 2396) => x"00", (0 + 2397) => x"00", (0 + 2398) => x"00", (0 + 2399) => x"00", (0 + 2400) => x"00", (0 + 2401) => x"00", (0 + 2402) => x"00", (0 + 2403) => x"00", (0 + 2404) => x"00", (0 + 2405) => x"00", (0 + 2406) => x"00", (0 + 2407) => x"00", (0 + 2408) => x"00", (0 + 2409) => x"00", (0 + 2410) => x"00", (0 + 2411) => x"00", (0 + 2412) => x"00", (0 + 2413) => x"00", (0 + 2414) => x"00", (0 + 2415) => x"00", (0 + 2416) => x"00", (0 + 2417) => x"00", (0 + 2418) => x"00", (0 + 2419) => x"00", (0 + 2420) => x"00", (0 + 2421) => x"00", (0 + 2422) => x"00", (0 + 2423) => x"00", (0 + 2424) => x"00", (0 + 2425) => x"00", (0 + 2426) => x"00", (0 + 2427) => x"00", (0 + 2428) => x"00", (0 + 2429) => x"00", (0 + 2430) => x"00", (0 + 2431) => x"00", (0 + 2432) => x"00", (0 + 2433) => x"00", (0 + 2434) => x"00", (0 + 2435) => x"00", (0 + 2436) => x"00", (0 + 2437) => x"00", (0 + 2438) => x"00", (0 + 2439) => x"00", (0 + 2440) => x"00", (0 + 2441) => x"00", (0 + 2442) => x"00", (0 + 2443) => x"00", (0 + 2444) => x"00", (0 + 2445) => x"00", (0 + 2446) => x"00", (0 + 2447) => x"00", (0 + 2448) => x"00", (0 + 2449) => x"00", (0 + 2450) => x"00", (0 + 2451) => x"00", (0 + 2452) => x"00", (0 + 2453) => x"00", (0 + 2454) => x"00", (0 + 2455) => x"00", (0 + 2456) => x"00", (0 + 2457) => x"00", (0 + 2458) => x"00", (0 + 2459) => x"00", (0 + 2460) => x"00", (0 + 2461) => x"00", (0 + 2462) => x"00", (0 + 2463) => x"00", (0 + 2464) => x"00", (0 + 2465) => x"00", (0 + 2466) => x"00", (0 + 2467) => x"00", (0 + 2468) => x"00", (0 + 2469) => x"00", (0 + 2470) => x"00", (0 + 2471) => x"00", (0 + 2472) => x"00", (0 + 2473) => x"00", (0 + 2474) => x"00", (0 + 2475) => x"00", (0 + 2476) => x"00", (0 + 2477) => x"00", (0 + 2478) => x"00", (0 + 2479) => x"00", (0 + 2480) => x"00", (0 + 2481) => x"00", (0 + 2482) => x"00", (0 + 2483) => x"00", (0 + 2484) => x"00", (0 + 2485) => x"00", (0 + 2486) => x"00", (0 + 2487) => x"00", (0 + 2488) => x"00", (0 + 2489) => x"00", (0 + 2490) => x"00", (0 + 2491) => x"00", (0 + 2492) => x"00", (0 + 2493) => x"00", (0 + 2494) => x"00", (0 + 2495) => x"00", (0 + 2496) => x"00", (0 + 2497) => x"00", (0 + 2498) => x"00", (0 + 2499) => x"00", (0 + 2500) => x"00", (0 + 2501) => x"00", (0 + 2502) => x"00", (0 + 2503) => x"00", (0 + 2504) => x"00", (0 + 2505) => x"00", (0 + 2506) => x"00", (0 + 2507) => x"00", (0 + 2508) => x"00", (0 + 2509) => x"00", (0 + 2510) => x"00", (0 + 2511) => x"00", (0 + 2512) => x"00", (0 + 2513) => x"00", (0 + 2514) => x"00", (0 + 2515) => x"00", (0 + 2516) => x"00", (0 + 2517) => x"00", (0 + 2518) => x"00", (0 + 2519) => x"00", (0 + 2520) => x"00", (0 + 2521) => x"00", (0 + 2522) => x"00", (0 + 2523) => x"00", (0 + 2524) => x"00", (0 + 2525) => x"00", (0 + 2526) => x"00", (0 + 2527) => x"00", (0 + 2528) => x"00", (0 + 2529) => x"00", (0 + 2530) => x"00", (0 + 2531) => x"00", (0 + 2532) => x"00", (0 + 2533) => x"00", (0 + 2534) => x"00", (0 + 2535) => x"00", (0 + 2536) => x"00", (0 + 2537) => x"00", (0 + 2538) => x"00", (0 + 2539) => x"00", (0 + 2540) => x"00", (0 + 2541) => x"00", (0 + 2542) => x"00", (0 + 2543) => x"00", (0 + 2544) => x"00", (0 + 2545) => x"00", (0 + 2546) => x"00", (0 + 2547) => x"00", (0 + 2548) => x"00", (0 + 2549) => x"00", (0 + 2550) => x"00", (0 + 2551) => x"00", (0 + 2552) => x"00", (0 + 2553) => x"00", (0 + 2554) => x"00", (0 + 2555) => x"00", (0 + 2556) => x"00", (0 + 2557) => x"00", (0 + 2558) => x"00", (0 + 2559) => x"00", (0 + 2560) => x"00", (0 + 2561) => x"00", (0 + 2562) => x"00", (0 + 2563) => x"00", (0 + 2564) => x"00", (0 + 2565) => x"00", (0 + 2566) => x"00", (0 + 2567) => x"00", (0 + 2568) => x"00", (0 + 2569) => x"00", (0 + 2570) => x"00", (0 + 2571) => x"00", (0 + 2572) => x"00", (0 + 2573) => x"00", (0 + 2574) => x"00", (0 + 2575) => x"00", (0 + 2576) => x"00", (0 + 2577) => x"00", (0 + 2578) => x"00", (0 + 2579) => x"00", (0 + 2580) => x"00", (0 + 2581) => x"00", (0 + 2582) => x"00", (0 + 2583) => x"00", (0 + 2584) => x"00", (0 + 2585) => x"00", (0 + 2586) => x"00", (0 + 2587) => x"00", (0 + 2588) => x"00", (0 + 2589) => x"00", (0 + 2590) => x"00", (0 + 2591) => x"00", (0 + 2592) => x"00", (0 + 2593) => x"00", (0 + 2594) => x"00", (0 + 2595) => x"00", (0 + 2596) => x"00", (0 + 2597) => x"00", (0 + 2598) => x"00", (0 + 2599) => x"00", (0 + 2600) => x"00", (0 + 2601) => x"00", (0 + 2602) => x"00", (0 + 2603) => x"00", (0 + 2604) => x"00", (0 + 2605) => x"00", (0 + 2606) => x"00", (0 + 2607) => x"00", (0 + 2608) => x"00", (0 + 2609) => x"00", (0 + 2610) => x"00", (0 + 2611) => x"00", (0 + 2612) => x"00", (0 + 2613) => x"00", (0 + 2614) => x"00", (0 + 2615) => x"00", (0 + 2616) => x"00", (0 + 2617) => x"00", (0 + 2618) => x"00", (0 + 2619) => x"00", (0 + 2620) => x"00", (0 + 2621) => x"00", (0 + 2622) => x"00", (0 + 2623) => x"00", (0 + 2624) => x"00", (0 + 2625) => x"00", (0 + 2626) => x"00", (0 + 2627) => x"00", (0 + 2628) => x"00", (0 + 2629) => x"00", (0 + 2630) => x"00", (0 + 2631) => x"00", (0 + 2632) => x"00", (0 + 2633) => x"00", (0 + 2634) => x"00", (0 + 2635) => x"00", (0 + 2636) => x"00", (0 + 2637) => x"00", (0 + 2638) => x"00", (0 + 2639) => x"00", (0 + 2640) => x"00", (0 + 2641) => x"00", (0 + 2642) => x"00", (0 + 2643) => x"00", (0 + 2644) => x"00", (0 + 2645) => x"00", (0 + 2646) => x"00", (0 + 2647) => x"00", (0 + 2648) => x"00", (0 + 2649) => x"00", (0 + 2650) => x"00", (0 + 2651) => x"00", (0 + 2652) => x"00", (0 + 2653) => x"00", (0 + 2654) => x"00", (0 + 2655) => x"00", (0 + 2656) => x"00", (0 + 2657) => x"00", (0 + 2658) => x"00", (0 + 2659) => x"00", (0 + 2660) => x"00", (0 + 2661) => x"00", (0 + 2662) => x"00", (0 + 2663) => x"00", (0 + 2664) => x"00", (0 + 2665) => x"00", (0 + 2666) => x"00", (0 + 2667) => x"00", (0 + 2668) => x"00", (0 + 2669) => x"00", (0 + 2670) => x"00", (0 + 2671) => x"00", (0 + 2672) => x"00", (0 + 2673) => x"00", (0 + 2674) => x"00", (0 + 2675) => x"00", (0 + 2676) => x"00", (0 + 2677) => x"00", (0 + 2678) => x"00", (0 + 2679) => x"00", (0 + 2680) => x"00", (0 + 2681) => x"00", (0 + 2682) => x"00", (0 + 2683) => x"00", (0 + 2684) => x"00", (0 + 2685) => x"00", (0 + 2686) => x"00", (0 + 2687) => x"00", (0 + 2688) => x"00", (0 + 2689) => x"00", (0 + 2690) => x"00", (0 + 2691) => x"00", (0 + 2692) => x"00", (0 + 2693) => x"00", (0 + 2694) => x"00", (0 + 2695) => x"00", (0 + 2696) => x"00", (0 + 2697) => x"00", (0 + 2698) => x"00", (0 + 2699) => x"00", (0 + 2700) => x"00", (0 + 2701) => x"00", (0 + 2702) => x"00", (0 + 2703) => x"00", (0 + 2704) => x"00", (0 + 2705) => x"00", (0 + 2706) => x"00", (0 + 2707) => x"00", (0 + 2708) => x"00", (0 + 2709) => x"00", (0 + 2710) => x"00", (0 + 2711) => x"00", (0 + 2712) => x"00", (0 + 2713) => x"00", (0 + 2714) => x"00", (0 + 2715) => x"00", (0 + 2716) => x"00", (0 + 2717) => x"00", (0 + 2718) => x"00", (0 + 2719) => x"00", (0 + 2720) => x"00", (0 + 2721) => x"00", (0 + 2722) => x"00", (0 + 2723) => x"00", (0 + 2724) => x"00", (0 + 2725) => x"00", (0 + 2726) => x"00", (0 + 2727) => x"00", (0 + 2728) => x"00", (0 + 2729) => x"00", (0 + 2730) => x"00", (0 + 2731) => x"00", (0 + 2732) => x"00", (0 + 2733) => x"00", (0 + 2734) => x"00", (0 + 2735) => x"00", (0 + 2736) => x"00", (0 + 2737) => x"00", (0 + 2738) => x"00", (0 + 2739) => x"00", (0 + 2740) => x"00", (0 + 2741) => x"00", (0 + 2742) => x"00", (0 + 2743) => x"00", (0 + 2744) => x"00", (0 + 2745) => x"00", (0 + 2746) => x"00", (0 + 2747) => x"00", (0 + 2748) => x"00", (0 + 2749) => x"00", (0 + 2750) => x"00", (0 + 2751) => x"00", (0 + 2752) => x"00", (0 + 2753) => x"00", (0 + 2754) => x"00", (0 + 2755) => x"00", (0 + 2756) => x"00", (0 + 2757) => x"00", (0 + 2758) => x"00", (0 + 2759) => x"00", (0 + 2760) => x"00", (0 + 2761) => x"00", (0 + 2762) => x"00", (0 + 2763) => x"00", (0 + 2764) => x"00", (0 + 2765) => x"00", (0 + 2766) => x"00", (0 + 2767) => x"00", (0 + 2768) => x"00", (0 + 2769) => x"00", (0 + 2770) => x"00", (0 + 2771) => x"00", (0 + 2772) => x"00", (0 + 2773) => x"00", (0 + 2774) => x"00", (0 + 2775) => x"00", (0 + 2776) => x"00", (0 + 2777) => x"00", (0 + 2778) => x"00", (0 + 2779) => x"00", (0 + 2780) => x"00", (0 + 2781) => x"00", (0 + 2782) => x"00", (0 + 2783) => x"00", (0 + 2784) => x"00", (0 + 2785) => x"00", (0 + 2786) => x"00", (0 + 2787) => x"00", (0 + 2788) => x"00", (0 + 2789) => x"00", (0 + 2790) => x"00", (0 + 2791) => x"00", (0 + 2792) => x"00", (0 + 2793) => x"00", (0 + 2794) => x"00", (0 + 2795) => x"00", (0 + 2796) => x"00", (0 + 2797) => x"00", (0 + 2798) => x"00", (0 + 2799) => x"00", (0 + 2800) => x"00", (0 + 2801) => x"00", (0 + 2802) => x"00", (0 + 2803) => x"00", (0 + 2804) => x"00", (0 + 2805) => x"00", (0 + 2806) => x"00", (0 + 2807) => x"00", (0 + 2808) => x"00", (0 + 2809) => x"00", (0 + 2810) => x"00", (0 + 2811) => x"00", (0 + 2812) => x"00", (0 + 2813) => x"00", (0 + 2814) => x"00", (0 + 2815) => x"00", (0 + 2816) => x"00", (0 + 2817) => x"00", (0 + 2818) => x"00", (0 + 2819) => x"00", (0 + 2820) => x"00", (0 + 2821) => x"00", (0 + 2822) => x"00", (0 + 2823) => x"00", (0 + 2824) => x"00", (0 + 2825) => x"00", (0 + 2826) => x"00", (0 + 2827) => x"00", (0 + 2828) => x"00", (0 + 2829) => x"00", (0 + 2830) => x"00", (0 + 2831) => x"00", (0 + 2832) => x"00", (0 + 2833) => x"00", (0 + 2834) => x"00", (0 + 2835) => x"00", (0 + 2836) => x"00", (0 + 2837) => x"00", (0 + 2838) => x"00", (0 + 2839) => x"00", (0 + 2840) => x"00", (0 + 2841) => x"00", (0 + 2842) => x"00", (0 + 2843) => x"00", (0 + 2844) => x"00", (0 + 2845) => x"00", (0 + 2846) => x"00", (0 + 2847) => x"00", (0 + 2848) => x"00", (0 + 2849) => x"00", (0 + 2850) => x"00", (0 + 2851) => x"00", (0 + 2852) => x"00", (0 + 2853) => x"00", (0 + 2854) => x"00", (0 + 2855) => x"00", (0 + 2856) => x"00", (0 + 2857) => x"00", (0 + 2858) => x"00", (0 + 2859) => x"00", (0 + 2860) => x"00", (0 + 2861) => x"00", (0 + 2862) => x"00", (0 + 2863) => x"00", (0 + 2864) => x"00", (0 + 2865) => x"00", (0 + 2866) => x"00", (0 + 2867) => x"00", (0 + 2868) => x"00", (0 + 2869) => x"00", (0 + 2870) => x"00", (0 + 2871) => x"00", (0 + 2872) => x"00", (0 + 2873) => x"00", (0 + 2874) => x"00", (0 + 2875) => x"00", (0 + 2876) => x"00", (0 + 2877) => x"00", (0 + 2878) => x"00", (0 + 2879) => x"00", (0 + 2880) => x"00", (0 + 2881) => x"00", (0 + 2882) => x"00", (0 + 2883) => x"00", (0 + 2884) => x"00", (0 + 2885) => x"00", (0 + 2886) => x"00", (0 + 2887) => x"00", (0 + 2888) => x"00", (0 + 2889) => x"00", (0 + 2890) => x"00", (0 + 2891) => x"00", (0 + 2892) => x"00", (0 + 2893) => x"00", (0 + 2894) => x"00", (0 + 2895) => x"00", (0 + 2896) => x"00", (0 + 2897) => x"00", (0 + 2898) => x"00", (0 + 2899) => x"00", (0 + 2900) => x"00", (0 + 2901) => x"00", (0 + 2902) => x"00", (0 + 2903) => x"00", (0 + 2904) => x"00", (0 + 2905) => x"00", (0 + 2906) => x"00", (0 + 2907) => x"00", (0 + 2908) => x"00", (0 + 2909) => x"00", (0 + 2910) => x"00", (0 + 2911) => x"00", (0 + 2912) => x"00", (0 + 2913) => x"00", (0 + 2914) => x"00", (0 + 2915) => x"00", (0 + 2916) => x"00", (0 + 2917) => x"00", (0 + 2918) => x"00", (0 + 2919) => x"00", (0 + 2920) => x"00", (0 + 2921) => x"00", (0 + 2922) => x"00", (0 + 2923) => x"00", (0 + 2924) => x"00", (0 + 2925) => x"00", (0 + 2926) => x"00", (0 + 2927) => x"00", (0 + 2928) => x"00", (0 + 2929) => x"00", (0 + 2930) => x"00", (0 + 2931) => x"00", (0 + 2932) => x"00", (0 + 2933) => x"00", (0 + 2934) => x"00", (0 + 2935) => x"00", (0 + 2936) => x"00", (0 + 2937) => x"00", (0 + 2938) => x"00", (0 + 2939) => x"00", (0 + 2940) => x"00", (0 + 2941) => x"00", (0 + 2942) => x"00", (0 + 2943) => x"00", (0 + 2944) => x"00", (0 + 2945) => x"00", (0 + 2946) => x"00", (0 + 2947) => x"00", (0 + 2948) => x"00", (0 + 2949) => x"00", (0 + 2950) => x"00", (0 + 2951) => x"00", (0 + 2952) => x"00", (0 + 2953) => x"00", (0 + 2954) => x"00", (0 + 2955) => x"00", (0 + 2956) => x"00", (0 + 2957) => x"00", (0 + 2958) => x"00", (0 + 2959) => x"00", (0 + 2960) => x"00", (0 + 2961) => x"00", (0 + 2962) => x"00", (0 + 2963) => x"00", (0 + 2964) => x"00", (0 + 2965) => x"00", (0 + 2966) => x"00", (0 + 2967) => x"00", (0 + 2968) => x"00", (0 + 2969) => x"00", (0 + 2970) => x"00", (0 + 2971) => x"00", (0 + 2972) => x"00", (0 + 2973) => x"00", (0 + 2974) => x"00", (0 + 2975) => x"00", (0 + 2976) => x"00", (0 + 2977) => x"00", (0 + 2978) => x"00", (0 + 2979) => x"00", (0 + 2980) => x"00", (0 + 2981) => x"00", (0 + 2982) => x"00", (0 + 2983) => x"00", (0 + 2984) => x"00", (0 + 2985) => x"00", (0 + 2986) => x"00", (0 + 2987) => x"00", (0 + 2988) => x"00", (0 + 2989) => x"00", (0 + 2990) => x"00", (0 + 2991) => x"00", (0 + 2992) => x"00", (0 + 2993) => x"00", (0 + 2994) => x"00", (0 + 2995) => x"00", (0 + 2996) => x"00", (0 + 2997) => x"00", (0 + 2998) => x"00", (0 + 2999) => x"00", (0 + 3000) => x"00", (0 + 3001) => x"00", (0 + 3002) => x"00", (0 + 3003) => x"00", (0 + 3004) => x"00", (0 + 3005) => x"00", (0 + 3006) => x"00", (0 + 3007) => x"00", (0 + 3008) => x"00", (0 + 3009) => x"00", (0 + 3010) => x"00", (0 + 3011) => x"00", (0 + 3012) => x"00", (0 + 3013) => x"00", (0 + 3014) => x"00", (0 + 3015) => x"00", (0 + 3016) => x"00", (0 + 3017) => x"00", (0 + 3018) => x"00", (0 + 3019) => x"00", (0 + 3020) => x"00", (0 + 3021) => x"00", (0 + 3022) => x"00", (0 + 3023) => x"00", (0 + 3024) => x"00", (0 + 3025) => x"00", (0 + 3026) => x"00", (0 + 3027) => x"00", (0 + 3028) => x"00", (0 + 3029) => x"00", (0 + 3030) => x"00", (0 + 3031) => x"00", (0 + 3032) => x"00", (0 + 3033) => x"00", (0 + 3034) => x"00", (0 + 3035) => x"00", (0 + 3036) => x"00", (0 + 3037) => x"00", (0 + 3038) => x"00", (0 + 3039) => x"00", (0 + 3040) => x"00", (0 + 3041) => x"00", (0 + 3042) => x"00", (0 + 3043) => x"00", (0 + 3044) => x"00", (0 + 3045) => x"00", (0 + 3046) => x"00", (0 + 3047) => x"00", (0 + 3048) => x"00", (0 + 3049) => x"00", (0 + 3050) => x"00", (0 + 3051) => x"00", (0 + 3052) => x"00", (0 + 3053) => x"00", (0 + 3054) => x"00", (0 + 3055) => x"00", (0 + 3056) => x"00", (0 + 3057) => x"00", (0 + 3058) => x"00", (0 + 3059) => x"00", (0 + 3060) => x"00", (0 + 3061) => x"00", (0 + 3062) => x"00", (0 + 3063) => x"00", (0 + 3064) => x"00", (0 + 3065) => x"00", (0 + 3066) => x"00", (0 + 3067) => x"00", (0 + 3068) => x"00", (0 + 3069) => x"00", (0 + 3070) => x"00", (0 + 3071) => x"00", (0 + 3072) => x"00", (0 + 3073) => x"00", (0 + 3074) => x"00", (0 + 3075) => x"00", (0 + 3076) => x"00", (0 + 3077) => x"00", (0 + 3078) => x"00", (0 + 3079) => x"00", (0 + 3080) => x"00", (0 + 3081) => x"00", (0 + 3082) => x"00", (0 + 3083) => x"00", (0 + 3084) => x"00", (0 + 3085) => x"00", (0 + 3086) => x"00", (0 + 3087) => x"00", (0 + 3088) => x"00", (0 + 3089) => x"00", (0 + 3090) => x"00", (0 + 3091) => x"00", (0 + 3092) => x"00", (0 + 3093) => x"00", (0 + 3094) => x"00", (0 + 3095) => x"00", (0 + 3096) => x"00", (0 + 3097) => x"00", (0 + 3098) => x"00", (0 + 3099) => x"00", (0 + 3100) => x"00", (0 + 3101) => x"00", (0 + 3102) => x"00", (0 + 3103) => x"00", (0 + 3104) => x"00", (0 + 3105) => x"00", (0 + 3106) => x"00", (0 + 3107) => x"00", (0 + 3108) => x"00", (0 + 3109) => x"00", (0 + 3110) => x"00", (0 + 3111) => x"00", (0 + 3112) => x"00", (0 + 3113) => x"00", (0 + 3114) => x"00", (0 + 3115) => x"00", (0 + 3116) => x"00", (0 + 3117) => x"00", (0 + 3118) => x"00", (0 + 3119) => x"00", (0 + 3120) => x"00", (0 + 3121) => x"00", (0 + 3122) => x"00", (0 + 3123) => x"00", (0 + 3124) => x"00", (0 + 3125) => x"00", (0 + 3126) => x"00", (0 + 3127) => x"00", (0 + 3128) => x"00", (0 + 3129) => x"00", (0 + 3130) => x"00", (0 + 3131) => x"00", (0 + 3132) => x"00", (0 + 3133) => x"00", (0 + 3134) => x"00", (0 + 3135) => x"00", (0 + 3136) => x"00", (0 + 3137) => x"00", (0 + 3138) => x"00", (0 + 3139) => x"00", (0 + 3140) => x"00", (0 + 3141) => x"00", (0 + 3142) => x"00", (0 + 3143) => x"00", (0 + 3144) => x"00", (0 + 3145) => x"00", (0 + 3146) => x"00", (0 + 3147) => x"00", (0 + 3148) => x"00", (0 + 3149) => x"00", (0 + 3150) => x"00", (0 + 3151) => x"00", (0 + 3152) => x"00", (0 + 3153) => x"00", (0 + 3154) => x"00", (0 + 3155) => x"00", (0 + 3156) => x"00", (0 + 3157) => x"00", (0 + 3158) => x"00", (0 + 3159) => x"00", (0 + 3160) => x"00", (0 + 3161) => x"00", (0 + 3162) => x"00", (0 + 3163) => x"00", (0 + 3164) => x"00", (0 + 3165) => x"00", (0 + 3166) => x"00", (0 + 3167) => x"00", (0 + 3168) => x"00", (0 + 3169) => x"00", (0 + 3170) => x"00", (0 + 3171) => x"00", (0 + 3172) => x"00", (0 + 3173) => x"00", (0 + 3174) => x"00", (0 + 3175) => x"00", (0 + 3176) => x"00", (0 + 3177) => x"00", (0 + 3178) => x"00", (0 + 3179) => x"00", (0 + 3180) => x"00", (0 + 3181) => x"00", (0 + 3182) => x"00", (0 + 3183) => x"00", (0 + 3184) => x"00", (0 + 3185) => x"00", (0 + 3186) => x"00", (0 + 3187) => x"00", (0 + 3188) => x"00", (0 + 3189) => x"00", (0 + 3190) => x"00", (0 + 3191) => x"00", (0 + 3192) => x"00", (0 + 3193) => x"00", (0 + 3194) => x"00", (0 + 3195) => x"00", (0 + 3196) => x"00", (0 + 3197) => x"00", (0 + 3198) => x"00", (0 + 3199) => x"00", (0 + 3200) => x"00", (0 + 3201) => x"00", (0 + 3202) => x"00", (0 + 3203) => x"00", (0 + 3204) => x"00", (0 + 3205) => x"00", (0 + 3206) => x"00", (0 + 3207) => x"00", (0 + 3208) => x"00", (0 + 3209) => x"00", (0 + 3210) => x"00", (0 + 3211) => x"00", (0 + 3212) => x"00", (0 + 3213) => x"00", (0 + 3214) => x"00", (0 + 3215) => x"00", (0 + 3216) => x"00", (0 + 3217) => x"00", (0 + 3218) => x"00", (0 + 3219) => x"00", (0 + 3220) => x"00", (0 + 3221) => x"00", (0 + 3222) => x"00", (0 + 3223) => x"00", (0 + 3224) => x"00", (0 + 3225) => x"00", (0 + 3226) => x"00", (0 + 3227) => x"00", (0 + 3228) => x"00", (0 + 3229) => x"00", (0 + 3230) => x"00", (0 + 3231) => x"00", (0 + 3232) => x"00", (0 + 3233) => x"00", (0 + 3234) => x"00", (0 + 3235) => x"00", (0 + 3236) => x"00", (0 + 3237) => x"00", (0 + 3238) => x"00", (0 + 3239) => x"00", (0 + 3240) => x"00", (0 + 3241) => x"00", (0 + 3242) => x"00", (0 + 3243) => x"00", (0 + 3244) => x"00", (0 + 3245) => x"00", (0 + 3246) => x"00", (0 + 3247) => x"00", (0 + 3248) => x"00", (0 + 3249) => x"00", (0 + 3250) => x"00", (0 + 3251) => x"00", (0 + 3252) => x"00", (0 + 3253) => x"00", (0 + 3254) => x"00", (0 + 3255) => x"00", (0 + 3256) => x"00", (0 + 3257) => x"00", (0 + 3258) => x"00", (0 + 3259) => x"00", (0 + 3260) => x"00", (0 + 3261) => x"00", (0 + 3262) => x"00", (0 + 3263) => x"00", (0 + 3264) => x"00", (0 + 3265) => x"00", (0 + 3266) => x"00", (0 + 3267) => x"00", (0 + 3268) => x"00", (0 + 3269) => x"00", (0 + 3270) => x"00", (0 + 3271) => x"00", (0 + 3272) => x"00", (0 + 3273) => x"00", (0 + 3274) => x"00", (0 + 3275) => x"00", (0 + 3276) => x"00", (0 + 3277) => x"00", (0 + 3278) => x"00", (0 + 3279) => x"00", (0 + 3280) => x"00", (0 + 3281) => x"00", (0 + 3282) => x"00", (0 + 3283) => x"00", (0 + 3284) => x"00", (0 + 3285) => x"00", (0 + 3286) => x"00", (0 + 3287) => x"00", (0 + 3288) => x"00", (0 + 3289) => x"00", (0 + 3290) => x"00", (0 + 3291) => x"00", (0 + 3292) => x"00", (0 + 3293) => x"00", (0 + 3294) => x"00", (0 + 3295) => x"00", (0 + 3296) => x"00", (0 + 3297) => x"00", (0 + 3298) => x"00", (0 + 3299) => x"00", (0 + 3300) => x"00", (0 + 3301) => x"00", (0 + 3302) => x"00", (0 + 3303) => x"00", (0 + 3304) => x"00", (0 + 3305) => x"00", (0 + 3306) => x"00", (0 + 3307) => x"00", (0 + 3308) => x"00", (0 + 3309) => x"00", (0 + 3310) => x"00", (0 + 3311) => x"00", (0 + 3312) => x"00", (0 + 3313) => x"00", (0 + 3314) => x"00", (0 + 3315) => x"00", (0 + 3316) => x"00", (0 + 3317) => x"00", (0 + 3318) => x"00", (0 + 3319) => x"00", (0 + 3320) => x"00", (0 + 3321) => x"00", (0 + 3322) => x"00", (0 + 3323) => x"00", (0 + 3324) => x"00", (0 + 3325) => x"00", (0 + 3326) => x"00", (0 + 3327) => x"00", (0 + 3328) => x"00", (0 + 3329) => x"00", (0 + 3330) => x"00", (0 + 3331) => x"00", (0 + 3332) => x"00", (0 + 3333) => x"00", (0 + 3334) => x"00", (0 + 3335) => x"00", (0 + 3336) => x"00", (0 + 3337) => x"00", (0 + 3338) => x"00", (0 + 3339) => x"00", (0 + 3340) => x"00", (0 + 3341) => x"00", (0 + 3342) => x"00", (0 + 3343) => x"00", (0 + 3344) => x"00", (0 + 3345) => x"00", (0 + 3346) => x"00", (0 + 3347) => x"00", (0 + 3348) => x"00", (0 + 3349) => x"00", (0 + 3350) => x"00", (0 + 3351) => x"00", (0 + 3352) => x"00", (0 + 3353) => x"00", (0 + 3354) => x"00", (0 + 3355) => x"00", (0 + 3356) => x"00", (0 + 3357) => x"00", (0 + 3358) => x"00", (0 + 3359) => x"00", (0 + 3360) => x"00", (0 + 3361) => x"00", (0 + 3362) => x"00", (0 + 3363) => x"00", (0 + 3364) => x"00", (0 + 3365) => x"00", (0 + 3366) => x"00", (0 + 3367) => x"00", (0 + 3368) => x"00", (0 + 3369) => x"00", (0 + 3370) => x"00", (0 + 3371) => x"00", (0 + 3372) => x"00", (0 + 3373) => x"00", (0 + 3374) => x"00", (0 + 3375) => x"00", (0 + 3376) => x"00", (0 + 3377) => x"00", (0 + 3378) => x"00", (0 + 3379) => x"00", (0 + 3380) => x"00", (0 + 3381) => x"00", (0 + 3382) => x"00", (0 + 3383) => x"00", (0 + 3384) => x"00", (0 + 3385) => x"00", (0 + 3386) => x"00", (0 + 3387) => x"00", (0 + 3388) => x"00", (0 + 3389) => x"00", (0 + 3390) => x"00", (0 + 3391) => x"00", (0 + 3392) => x"00", (0 + 3393) => x"00", (0 + 3394) => x"00", (0 + 3395) => x"00", (0 + 3396) => x"00", (0 + 3397) => x"00", (0 + 3398) => x"00", (0 + 3399) => x"00", (0 + 3400) => x"00", (0 + 3401) => x"00", (0 + 3402) => x"00", (0 + 3403) => x"00", (0 + 3404) => x"00", (0 + 3405) => x"00", (0 + 3406) => x"00", (0 + 3407) => x"00", (0 + 3408) => x"00", (0 + 3409) => x"00", (0 + 3410) => x"00", (0 + 3411) => x"00", (0 + 3412) => x"00", (0 + 3413) => x"00", (0 + 3414) => x"00", (0 + 3415) => x"00", (0 + 3416) => x"00", (0 + 3417) => x"00", (0 + 3418) => x"00", (0 + 3419) => x"00", (0 + 3420) => x"00", (0 + 3421) => x"00", (0 + 3422) => x"00", (0 + 3423) => x"00", (0 + 3424) => x"00", (0 + 3425) => x"00", (0 + 3426) => x"00", (0 + 3427) => x"00", (0 + 3428) => x"00", (0 + 3429) => x"00", (0 + 3430) => x"00", (0 + 3431) => x"00", (0 + 3432) => x"00", (0 + 3433) => x"00", (0 + 3434) => x"00", (0 + 3435) => x"00", (0 + 3436) => x"00", (0 + 3437) => x"00", (0 + 3438) => x"00", (0 + 3439) => x"00", (0 + 3440) => x"00", (0 + 3441) => x"00", (0 + 3442) => x"00", (0 + 3443) => x"00", (0 + 3444) => x"00", (0 + 3445) => x"00", (0 + 3446) => x"00", (0 + 3447) => x"00", (0 + 3448) => x"00", (0 + 3449) => x"00", (0 + 3450) => x"00", (0 + 3451) => x"00", (0 + 3452) => x"00", (0 + 3453) => x"00", (0 + 3454) => x"00", (0 + 3455) => x"00", (0 + 3456) => x"00", (0 + 3457) => x"00", (0 + 3458) => x"00", (0 + 3459) => x"00", (0 + 3460) => x"00", (0 + 3461) => x"00", (0 + 3462) => x"00", (0 + 3463) => x"00", (0 + 3464) => x"00", (0 + 3465) => x"00", (0 + 3466) => x"00", (0 + 3467) => x"00", (0 + 3468) => x"00", (0 + 3469) => x"00", (0 + 3470) => x"00", (0 + 3471) => x"00", (0 + 3472) => x"00", (0 + 3473) => x"00", (0 + 3474) => x"00", (0 + 3475) => x"00", (0 + 3476) => x"00", (0 + 3477) => x"00", (0 + 3478) => x"00", (0 + 3479) => x"00", (0 + 3480) => x"00", (0 + 3481) => x"00", (0 + 3482) => x"00", (0 + 3483) => x"00", (0 + 3484) => x"00", (0 + 3485) => x"00", (0 + 3486) => x"00", (0 + 3487) => x"00", (0 + 3488) => x"00", (0 + 3489) => x"00", (0 + 3490) => x"00", (0 + 3491) => x"00", (0 + 3492) => x"00", (0 + 3493) => x"00", (0 + 3494) => x"00", (0 + 3495) => x"00", (0 + 3496) => x"00", (0 + 3497) => x"00", (0 + 3498) => x"00", (0 + 3499) => x"00", (0 + 3500) => x"00", (0 + 3501) => x"00", (0 + 3502) => x"00", (0 + 3503) => x"00", (0 + 3504) => x"00", (0 + 3505) => x"00", (0 + 3506) => x"00", (0 + 3507) => x"00", (0 + 3508) => x"00", (0 + 3509) => x"00", (0 + 3510) => x"00", (0 + 3511) => x"00", (0 + 3512) => x"00", (0 + 3513) => x"00", (0 + 3514) => x"00", (0 + 3515) => x"00", (0 + 3516) => x"00", (0 + 3517) => x"00", (0 + 3518) => x"00", (0 + 3519) => x"00", (0 + 3520) => x"00", (0 + 3521) => x"00", (0 + 3522) => x"00", (0 + 3523) => x"00", (0 + 3524) => x"00", (0 + 3525) => x"00", (0 + 3526) => x"00", (0 + 3527) => x"00", (0 + 3528) => x"00", (0 + 3529) => x"00", (0 + 3530) => x"00", (0 + 3531) => x"00", (0 + 3532) => x"00", (0 + 3533) => x"00", (0 + 3534) => x"00", (0 + 3535) => x"00", (0 + 3536) => x"00", (0 + 3537) => x"00", (0 + 3538) => x"00", (0 + 3539) => x"00", (0 + 3540) => x"00", (0 + 3541) => x"00", (0 + 3542) => x"00", (0 + 3543) => x"00", (0 + 3544) => x"00", (0 + 3545) => x"00", (0 + 3546) => x"00", (0 + 3547) => x"00", (0 + 3548) => x"00", (0 + 3549) => x"00", (0 + 3550) => x"00", (0 + 3551) => x"00", (0 + 3552) => x"00", (0 + 3553) => x"00", (0 + 3554) => x"00", (0 + 3555) => x"00", (0 + 3556) => x"00", (0 + 3557) => x"00", (0 + 3558) => x"00", (0 + 3559) => x"00", (0 + 3560) => x"00", (0 + 3561) => x"00", (0 + 3562) => x"00", (0 + 3563) => x"00", (0 + 3564) => x"00", (0 + 3565) => x"00", (0 + 3566) => x"00", (0 + 3567) => x"00", (0 + 3568) => x"00", (0 + 3569) => x"00", (0 + 3570) => x"00", (0 + 3571) => x"00", (0 + 3572) => x"00", (0 + 3573) => x"00", (0 + 3574) => x"00", (0 + 3575) => x"00", (0 + 3576) => x"00", (0 + 3577) => x"00", (0 + 3578) => x"00", (0 + 3579) => x"00", (0 + 3580) => x"00", (0 + 3581) => x"00", (0 + 3582) => x"00", (0 + 3583) => x"00", (0 + 3584) => x"00", (0 + 3585) => x"00", (0 + 3586) => x"00", (0 + 3587) => x"00", (0 + 3588) => x"00", (0 + 3589) => x"00", (0 + 3590) => x"00", (0 + 3591) => x"00", (0 + 3592) => x"00", (0 + 3593) => x"00", (0 + 3594) => x"00", (0 + 3595) => x"00", (0 + 3596) => x"00", (0 + 3597) => x"00", (0 + 3598) => x"00", (0 + 3599) => x"00", (0 + 3600) => x"00", (0 + 3601) => x"00", (0 + 3602) => x"00", (0 + 3603) => x"00", (0 + 3604) => x"00", (0 + 3605) => x"00", (0 + 3606) => x"00", (0 + 3607) => x"00", (0 + 3608) => x"00", (0 + 3609) => x"00", (0 + 3610) => x"00", (0 + 3611) => x"00", (0 + 3612) => x"00", (0 + 3613) => x"00", (0 + 3614) => x"00", (0 + 3615) => x"00", (0 + 3616) => x"00", (0 + 3617) => x"00", (0 + 3618) => x"00", (0 + 3619) => x"00", (0 + 3620) => x"00", (0 + 3621) => x"00", (0 + 3622) => x"00", (0 + 3623) => x"00", (0 + 3624) => x"00", (0 + 3625) => x"00", (0 + 3626) => x"00", (0 + 3627) => x"00", (0 + 3628) => x"00", (0 + 3629) => x"00", (0 + 3630) => x"00", (0 + 3631) => x"00", (0 + 3632) => x"00", (0 + 3633) => x"00", (0 + 3634) => x"00", (0 + 3635) => x"00", (0 + 3636) => x"00", (0 + 3637) => x"00", (0 + 3638) => x"00", (0 + 3639) => x"00", (0 + 3640) => x"00", (0 + 3641) => x"00", (0 + 3642) => x"00", (0 + 3643) => x"00", (0 + 3644) => x"00", (0 + 3645) => x"00", (0 + 3646) => x"00", (0 + 3647) => x"00", (0 + 3648) => x"00", (0 + 3649) => x"00", (0 + 3650) => x"00", (0 + 3651) => x"00", (0 + 3652) => x"00", (0 + 3653) => x"00", (0 + 3654) => x"00", (0 + 3655) => x"00", (0 + 3656) => x"00", (0 + 3657) => x"00", (0 + 3658) => x"00", (0 + 3659) => x"00", (0 + 3660) => x"00", (0 + 3661) => x"00", (0 + 3662) => x"00", (0 + 3663) => x"00", (0 + 3664) => x"00", (0 + 3665) => x"00", (0 + 3666) => x"00", (0 + 3667) => x"00", (0 + 3668) => x"00", (0 + 3669) => x"00", (0 + 3670) => x"00", (0 + 3671) => x"00", (0 + 3672) => x"00", (0 + 3673) => x"00", (0 + 3674) => x"00", (0 + 3675) => x"00", (0 + 3676) => x"00", (0 + 3677) => x"00", (0 + 3678) => x"00", (0 + 3679) => x"00", (0 + 3680) => x"00", (0 + 3681) => x"00", (0 + 3682) => x"00", (0 + 3683) => x"00", (0 + 3684) => x"00", (0 + 3685) => x"00", (0 + 3686) => x"00", (0 + 3687) => x"00", (0 + 3688) => x"00", (0 + 3689) => x"00", (0 + 3690) => x"00", (0 + 3691) => x"00", (0 + 3692) => x"00", (0 + 3693) => x"00", (0 + 3694) => x"00", (0 + 3695) => x"00", (0 + 3696) => x"00", (0 + 3697) => x"00", (0 + 3698) => x"00", (0 + 3699) => x"00", (0 + 3700) => x"00", (0 + 3701) => x"00", (0 + 3702) => x"00", (0 + 3703) => x"00", (0 + 3704) => x"00", (0 + 3705) => x"00", (0 + 3706) => x"00", (0 + 3707) => x"00", (0 + 3708) => x"00", (0 + 3709) => x"00", (0 + 3710) => x"00", (0 + 3711) => x"00", (0 + 3712) => x"00", (0 + 3713) => x"00", (0 + 3714) => x"00", (0 + 3715) => x"00", (0 + 3716) => x"00", (0 + 3717) => x"00", (0 + 3718) => x"00", (0 + 3719) => x"00", (0 + 3720) => x"00", (0 + 3721) => x"00", (0 + 3722) => x"00", (0 + 3723) => x"00", (0 + 3724) => x"00", (0 + 3725) => x"00", (0 + 3726) => x"00", (0 + 3727) => x"00", (0 + 3728) => x"00", (0 + 3729) => x"00", (0 + 3730) => x"00", (0 + 3731) => x"00", (0 + 3732) => x"00", (0 + 3733) => x"00", (0 + 3734) => x"00", (0 + 3735) => x"00", (0 + 3736) => x"00", (0 + 3737) => x"00", (0 + 3738) => x"00", (0 + 3739) => x"00", (0 + 3740) => x"00", (0 + 3741) => x"00", (0 + 3742) => x"00", (0 + 3743) => x"00", (0 + 3744) => x"00", (0 + 3745) => x"00", (0 + 3746) => x"00", (0 + 3747) => x"00", (0 + 3748) => x"00", (0 + 3749) => x"00", (0 + 3750) => x"00", (0 + 3751) => x"00", (0 + 3752) => x"00", (0 + 3753) => x"00", (0 + 3754) => x"00", (0 + 3755) => x"00", (0 + 3756) => x"00", (0 + 3757) => x"00", (0 + 3758) => x"00", (0 + 3759) => x"00", (0 + 3760) => x"00", (0 + 3761) => x"00", (0 + 3762) => x"00", (0 + 3763) => x"00", (0 + 3764) => x"00", (0 + 3765) => x"00", (0 + 3766) => x"00", (0 + 3767) => x"00", (0 + 3768) => x"00", (0 + 3769) => x"00", (0 + 3770) => x"00", (0 + 3771) => x"00", (0 + 3772) => x"00", (0 + 3773) => x"00", (0 + 3774) => x"00", (0 + 3775) => x"00", (0 + 3776) => x"00", (0 + 3777) => x"00", (0 + 3778) => x"00", (0 + 3779) => x"00", (0 + 3780) => x"00", (0 + 3781) => x"00", (0 + 3782) => x"00", (0 + 3783) => x"00", (0 + 3784) => x"00", (0 + 3785) => x"00", (0 + 3786) => x"00", (0 + 3787) => x"00", (0 + 3788) => x"00", (0 + 3789) => x"00", (0 + 3790) => x"00", (0 + 3791) => x"00", (0 + 3792) => x"00", (0 + 3793) => x"00", (0 + 3794) => x"00", (0 + 3795) => x"00", (0 + 3796) => x"00", (0 + 3797) => x"00", (0 + 3798) => x"00", (0 + 3799) => x"00", (0 + 3800) => x"00", (0 + 3801) => x"00", (0 + 3802) => x"00", (0 + 3803) => x"00", (0 + 3804) => x"00", (0 + 3805) => x"00", (0 + 3806) => x"00", (0 + 3807) => x"00", (0 + 3808) => x"00", (0 + 3809) => x"00", (0 + 3810) => x"00", (0 + 3811) => x"00", (0 + 3812) => x"00", (0 + 3813) => x"00", (0 + 3814) => x"00", (0 + 3815) => x"00", (0 + 3816) => x"00", (0 + 3817) => x"00", (0 + 3818) => x"00", (0 + 3819) => x"00", (0 + 3820) => x"00", (0 + 3821) => x"00", (0 + 3822) => x"00", (0 + 3823) => x"00", (0 + 3824) => x"00", (0 + 3825) => x"00", (0 + 3826) => x"00", (0 + 3827) => x"00", (0 + 3828) => x"00", (0 + 3829) => x"00", (0 + 3830) => x"00", (0 + 3831) => x"00", (0 + 3832) => x"00", (0 + 3833) => x"00", (0 + 3834) => x"00", (0 + 3835) => x"00", (0 + 3836) => x"00", (0 + 3837) => x"00", (0 + 3838) => x"00", (0 + 3839) => x"00", (0 + 3840) => x"00", (0 + 3841) => x"00", (0 + 3842) => x"00", (0 + 3843) => x"00", (0 + 3844) => x"00", (0 + 3845) => x"00", (0 + 3846) => x"00", (0 + 3847) => x"00", (0 + 3848) => x"00", (0 + 3849) => x"00", (0 + 3850) => x"00", (0 + 3851) => x"00", (0 + 3852) => x"00", (0 + 3853) => x"00", (0 + 3854) => x"00", (0 + 3855) => x"00", (0 + 3856) => x"00", (0 + 3857) => x"00", (0 + 3858) => x"00", (0 + 3859) => x"00", (0 + 3860) => x"00", (0 + 3861) => x"00", (0 + 3862) => x"00", (0 + 3863) => x"00", (0 + 3864) => x"00", (0 + 3865) => x"00", (0 + 3866) => x"00", (0 + 3867) => x"00", (0 + 3868) => x"00", (0 + 3869) => x"00", (0 + 3870) => x"00", (0 + 3871) => x"00", (0 + 3872) => x"00", (0 + 3873) => x"00", (0 + 3874) => x"00", (0 + 3875) => x"00", (0 + 3876) => x"00", (0 + 3877) => x"00", (0 + 3878) => x"00", (0 + 3879) => x"00", (0 + 3880) => x"00", (0 + 3881) => x"00", (0 + 3882) => x"00", (0 + 3883) => x"00", (0 + 3884) => x"00", (0 + 3885) => x"00", (0 + 3886) => x"00", (0 + 3887) => x"00", (0 + 3888) => x"00", (0 + 3889) => x"00", (0 + 3890) => x"00", (0 + 3891) => x"00", (0 + 3892) => x"00", (0 + 3893) => x"00", (0 + 3894) => x"00", (0 + 3895) => x"00", (0 + 3896) => x"00", (0 + 3897) => x"00", (0 + 3898) => x"00", (0 + 3899) => x"00", (0 + 3900) => x"00", (0 + 3901) => x"00", (0 + 3902) => x"00", (0 + 3903) => x"00", (0 + 3904) => x"00", (0 + 3905) => x"00", (0 + 3906) => x"00", (0 + 3907) => x"00", (0 + 3908) => x"00", (0 + 3909) => x"00", (0 + 3910) => x"00", (0 + 3911) => x"00", (0 + 3912) => x"00", (0 + 3913) => x"00", (0 + 3914) => x"00", (0 + 3915) => x"00", (0 + 3916) => x"00", (0 + 3917) => x"00", (0 + 3918) => x"00", (0 + 3919) => x"00", (0 + 3920) => x"00", (0 + 3921) => x"00", (0 + 3922) => x"00", (0 + 3923) => x"00", (0 + 3924) => x"00", (0 + 3925) => x"00", (0 + 3926) => x"00", (0 + 3927) => x"00", (0 + 3928) => x"00", (0 + 3929) => x"00", (0 + 3930) => x"00", (0 + 3931) => x"00", (0 + 3932) => x"00", (0 + 3933) => x"00", (0 + 3934) => x"00", (0 + 3935) => x"00", (0 + 3936) => x"00", (0 + 3937) => x"00", (0 + 3938) => x"00", (0 + 3939) => x"00", (0 + 3940) => x"00", (0 + 3941) => x"00", (0 + 3942) => x"00", (0 + 3943) => x"00", (0 + 3944) => x"00", (0 + 3945) => x"00", (0 + 3946) => x"00", (0 + 3947) => x"00", (0 + 3948) => x"00", (0 + 3949) => x"00", (0 + 3950) => x"00", (0 + 3951) => x"00", (0 + 3952) => x"00", (0 + 3953) => x"00", (0 + 3954) => x"00", (0 + 3955) => x"00", (0 + 3956) => x"00", (0 + 3957) => x"00", (0 + 3958) => x"00", (0 + 3959) => x"00", (0 + 3960) => x"00", (0 + 3961) => x"00", (0 + 3962) => x"00", (0 + 3963) => x"00", (0 + 3964) => x"00", (0 + 3965) => x"00", (0 + 3966) => x"00", (0 + 3967) => x"00", (0 + 3968) => x"00", (0 + 3969) => x"00", (0 + 3970) => x"00", (0 + 3971) => x"00", (0 + 3972) => x"00", (0 + 3973) => x"00", (0 + 3974) => x"00", (0 + 3975) => x"00", (0 + 3976) => x"00", (0 + 3977) => x"00", (0 + 3978) => x"00", (0 + 3979) => x"00", (0 + 3980) => x"00", (0 + 3981) => x"00", (0 + 3982) => x"00", (0 + 3983) => x"00", (0 + 3984) => x"00", (0 + 3985) => x"00", (0 + 3986) => x"00", (0 + 3987) => x"00", (0 + 3988) => x"00", (0 + 3989) => x"00", (0 + 3990) => x"00", (0 + 3991) => x"00", (0 + 3992) => x"00", (0 + 3993) => x"00", (0 + 3994) => x"00", (0 + 3995) => x"00", (0 + 3996) => x"00", (0 + 3997) => x"00", (0 + 3998) => x"00", (0 + 3999) => x"00", (0 + 4000) => x"00", (0 + 4001) => x"00", (0 + 4002) => x"00", (0 + 4003) => x"00", (0 + 4004) => x"00", (0 + 4005) => x"00", (0 + 4006) => x"00", (0 + 4007) => x"00", (0 + 4008) => x"00", (0 + 4009) => x"00", (0 + 4010) => x"00", (0 + 4011) => x"00", (0 + 4012) => x"00", (0 + 4013) => x"00", (0 + 4014) => x"00", (0 + 4015) => x"00", (0 + 4016) => x"00", (0 + 4017) => x"00", (0 + 4018) => x"00", (0 + 4019) => x"00", (0 + 4020) => x"00", (0 + 4021) => x"00", (0 + 4022) => x"00", (0 + 4023) => x"00", (0 + 4024) => x"00", (0 + 4025) => x"00", (0 + 4026) => x"00", (0 + 4027) => x"00", (0 + 4028) => x"00", (0 + 4029) => x"00", (0 + 4030) => x"00", (0 + 4031) => x"00", (0 + 4032) => x"00", (0 + 4033) => x"00", (0 + 4034) => x"00", (0 + 4035) => x"00", (0 + 4036) => x"00", (0 + 4037) => x"00", (0 + 4038) => x"00", (0 + 4039) => x"00", (0 + 4040) => x"00", (0 + 4041) => x"00", (0 + 4042) => x"00", (0 + 4043) => x"00", (0 + 4044) => x"00", (0 + 4045) => x"00", (0 + 4046) => x"00", (0 + 4047) => x"00", (0 + 4048) => x"00", (0 + 4049) => x"00", (0 + 4050) => x"00", (0 + 4051) => x"00", (0 + 4052) => x"00", (0 + 4053) => x"00", (0 + 4054) => x"00", (0 + 4055) => x"00", (0 + 4056) => x"00", (0 + 4057) => x"00", (0 + 4058) => x"00", (0 + 4059) => x"00", (0 + 4060) => x"00", (0 + 4061) => x"00", (0 + 4062) => x"00", (0 + 4063) => x"00", (0 + 4064) => x"00", (0 + 4065) => x"00", (0 + 4066) => x"00", (0 + 4067) => x"00", (0 + 4068) => x"00", (0 + 4069) => x"00", (0 + 4070) => x"00", (0 + 4071) => x"00", (0 + 4072) => x"00", (0 + 4073) => x"00", (0 + 4074) => x"00", (0 + 4075) => x"00", (0 + 4076) => x"00", (0 + 4077) => x"00", (0 + 4078) => x"00", (0 + 4079) => x"00", (0 + 4080) => x"00", (0 + 4081) => x"00", (0 + 4082) => x"00", (0 + 4083) => x"00", (0 + 4084) => x"00", (0 + 4085) => x"00", (0 + 4086) => x"00", (0 + 4087) => x"00", (0 + 4088) => x"00", (0 + 4089) => x"00", (0 + 4090) => x"00", (0 + 4091) => x"00", (0 + 4092) => x"00", (0 + 4093) => x"00", (0 + 4094) => x"00", (0 + 4095) => x"00", (0 + 4096) => x"00", (0 + 4097) => x"00", (0 + 4098) => x"00", (0 + 4099) => x"00", (0 + 4100) => x"00", (0 + 4101) => x"00", (0 + 4102) => x"00", (0 + 4103) => x"00", (0 + 4104) => x"00", (0 + 4105) => x"00", (0 + 4106) => x"00", (0 + 4107) => x"00", (0 + 4108) => x"00", (0 + 4109) => x"00", (0 + 4110) => x"00", (0 + 4111) => x"00", (0 + 4112) => x"00", (0 + 4113) => x"00", (0 + 4114) => x"00", (0 + 4115) => x"00", (0 + 4116) => x"00", (0 + 4117) => x"00", (0 + 4118) => x"00", (0 + 4119) => x"00", (0 + 4120) => x"00", (0 + 4121) => x"00", (0 + 4122) => x"00", (0 + 4123) => x"00", (0 + 4124) => x"00", (0 + 4125) => x"00", (0 + 4126) => x"00", (0 + 4127) => x"00", (0 + 4128) => x"00", (0 + 4129) => x"00", (0 + 4130) => x"00", (0 + 4131) => x"00", (0 + 4132) => x"00", (0 + 4133) => x"00", (0 + 4134) => x"00", (0 + 4135) => x"00", (0 + 4136) => x"00", (0 + 4137) => x"00", (0 + 4138) => x"00", (0 + 4139) => x"00", (0 + 4140) => x"00", (0 + 4141) => x"00", (0 + 4142) => x"00", (0 + 4143) => x"00", (0 + 4144) => x"00", (0 + 4145) => x"00", (0 + 4146) => x"00", (0 + 4147) => x"00", (0 + 4148) => x"00", (0 + 4149) => x"00", (0 + 4150) => x"00", (0 + 4151) => x"00", (0 + 4152) => x"00", (0 + 4153) => x"00", (0 + 4154) => x"00", (0 + 4155) => x"00", (0 + 4156) => x"00", (0 + 4157) => x"00", (0 + 4158) => x"00", (0 + 4159) => x"00", (0 + 4160) => x"00", (0 + 4161) => x"00", (0 + 4162) => x"00", (0 + 4163) => x"00", (0 + 4164) => x"00", (0 + 4165) => x"00", (0 + 4166) => x"00", (0 + 4167) => x"00", (0 + 4168) => x"00", (0 + 4169) => x"00", (0 + 4170) => x"00", (0 + 4171) => x"00", (0 + 4172) => x"00", (0 + 4173) => x"00", (0 + 4174) => x"00", (0 + 4175) => x"00", (0 + 4176) => x"00", (0 + 4177) => x"00", (0 + 4178) => x"00", (0 + 4179) => x"00", (0 + 4180) => x"00", (0 + 4181) => x"00", (0 + 4182) => x"00", (0 + 4183) => x"00", (0 + 4184) => x"00", (0 + 4185) => x"00", (0 + 4186) => x"00", (0 + 4187) => x"00", (0 + 4188) => x"00", (0 + 4189) => x"00", (0 + 4190) => x"00", (0 + 4191) => x"00", (0 + 4192) => x"00", (0 + 4193) => x"00", (0 + 4194) => x"00", (0 + 4195) => x"00", (0 + 4196) => x"00", (0 + 4197) => x"00", (0 + 4198) => x"00", (0 + 4199) => x"00", (0 + 4200) => x"00", (0 + 4201) => x"00", (0 + 4202) => x"00", (0 + 4203) => x"00", (0 + 4204) => x"00", (0 + 4205) => x"00", (0 + 4206) => x"00", (0 + 4207) => x"00", (0 + 4208) => x"00", (0 + 4209) => x"00", (0 + 4210) => x"00", (0 + 4211) => x"00", (0 + 4212) => x"00", (0 + 4213) => x"00", (0 + 4214) => x"00", (0 + 4215) => x"00", (0 + 4216) => x"00", (0 + 4217) => x"00", (0 + 4218) => x"00", (0 + 4219) => x"00", (0 + 4220) => x"00", (0 + 4221) => x"00", (0 + 4222) => x"00", (0 + 4223) => x"00", (0 + 4224) => x"00", (0 + 4225) => x"00", (0 + 4226) => x"00", (0 + 4227) => x"00", (0 + 4228) => x"00", (0 + 4229) => x"00", (0 + 4230) => x"00", (0 + 4231) => x"00", (0 + 4232) => x"00", (0 + 4233) => x"00", (0 + 4234) => x"00", (0 + 4235) => x"00", (0 + 4236) => x"00", (0 + 4237) => x"00", (0 + 4238) => x"00", (0 + 4239) => x"00", (0 + 4240) => x"00", (0 + 4241) => x"00", (0 + 4242) => x"00", (0 + 4243) => x"00", (0 + 4244) => x"00", (0 + 4245) => x"00", (0 + 4246) => x"00", (0 + 4247) => x"00", (0 + 4248) => x"00", (0 + 4249) => x"00", (0 + 4250) => x"00", (0 + 4251) => x"00", (0 + 4252) => x"00", (0 + 4253) => x"00", (0 + 4254) => x"00", (0 + 4255) => x"00", (0 + 4256) => x"00", (0 + 4257) => x"00", (0 + 4258) => x"00", (0 + 4259) => x"00", (0 + 4260) => x"00", (0 + 4261) => x"00", (0 + 4262) => x"00", (0 + 4263) => x"00", (0 + 4264) => x"00", (0 + 4265) => x"00", (0 + 4266) => x"00", (0 + 4267) => x"00", (0 + 4268) => x"00", (0 + 4269) => x"00", (0 + 4270) => x"00", (0 + 4271) => x"00", (0 + 4272) => x"00", (0 + 4273) => x"00", (0 + 4274) => x"00", (0 + 4275) => x"00", (0 + 4276) => x"00", (0 + 4277) => x"00", (0 + 4278) => x"00", (0 + 4279) => x"00", (0 + 4280) => x"00", (0 + 4281) => x"00", (0 + 4282) => x"00", (0 + 4283) => x"00", (0 + 4284) => x"00", (0 + 4285) => x"00", (0 + 4286) => x"00", (0 + 4287) => x"00", (0 + 4288) => x"00", (0 + 4289) => x"00", (0 + 4290) => x"00", (0 + 4291) => x"00", (0 + 4292) => x"00", (0 + 4293) => x"00", (0 + 4294) => x"00", (0 + 4295) => x"00", (0 + 4296) => x"00", (0 + 4297) => x"00", (0 + 4298) => x"00", (0 + 4299) => x"00", (0 + 4300) => x"00", (0 + 4301) => x"00", (0 + 4302) => x"00", (0 + 4303) => x"00", (0 + 4304) => x"00", (0 + 4305) => x"00", (0 + 4306) => x"00", (0 + 4307) => x"00", (0 + 4308) => x"00", (0 + 4309) => x"00", (0 + 4310) => x"00", (0 + 4311) => x"00", (0 + 4312) => x"00", (0 + 4313) => x"00", (0 + 4314) => x"00", (0 + 4315) => x"00", (0 + 4316) => x"00", (0 + 4317) => x"00", (0 + 4318) => x"00", (0 + 4319) => x"00", (0 + 4320) => x"00", (0 + 4321) => x"00", (0 + 4322) => x"00", (0 + 4323) => x"00", (0 + 4324) => x"00", (0 + 4325) => x"00", (0 + 4326) => x"00", (0 + 4327) => x"00", (0 + 4328) => x"00", (0 + 4329) => x"00", (0 + 4330) => x"00", (0 + 4331) => x"00", (0 + 4332) => x"00", (0 + 4333) => x"00", (0 + 4334) => x"00", (0 + 4335) => x"00", (0 + 4336) => x"00", (0 + 4337) => x"00", (0 + 4338) => x"00", (0 + 4339) => x"00", (0 + 4340) => x"00", (0 + 4341) => x"00", (0 + 4342) => x"00", (0 + 4343) => x"00", (0 + 4344) => x"00", (0 + 4345) => x"00", (0 + 4346) => x"00", (0 + 4347) => x"00", (0 + 4348) => x"00", (0 + 4349) => x"00", (0 + 4350) => x"00", (0 + 4351) => x"00", (0 + 4352) => x"00", (0 + 4353) => x"00", (0 + 4354) => x"00", (0 + 4355) => x"00", (0 + 4356) => x"00", (0 + 4357) => x"00", (0 + 4358) => x"00", (0 + 4359) => x"00", (0 + 4360) => x"00", (0 + 4361) => x"00", (0 + 4362) => x"00", (0 + 4363) => x"00", (0 + 4364) => x"00", (0 + 4365) => x"00", (0 + 4366) => x"00", (0 + 4367) => x"00", (0 + 4368) => x"00", (0 + 4369) => x"00", (0 + 4370) => x"00", (0 + 4371) => x"00", (0 + 4372) => x"00", (0 + 4373) => x"00", (0 + 4374) => x"00", (0 + 4375) => x"00", (0 + 4376) => x"00", (0 + 4377) => x"00", (0 + 4378) => x"00", (0 + 4379) => x"00", (0 + 4380) => x"00", (0 + 4381) => x"00", (0 + 4382) => x"00", (0 + 4383) => x"00", (0 + 4384) => x"00", (0 + 4385) => x"00", (0 + 4386) => x"00", (0 + 4387) => x"00", (0 + 4388) => x"00", (0 + 4389) => x"00", (0 + 4390) => x"00", (0 + 4391) => x"00", (0 + 4392) => x"00", (0 + 4393) => x"00", (0 + 4394) => x"00", (0 + 4395) => x"00", (0 + 4396) => x"00", (0 + 4397) => x"00", (0 + 4398) => x"00", (0 + 4399) => x"00", (0 + 4400) => x"00", (0 + 4401) => x"00", (0 + 4402) => x"00", (0 + 4403) => x"00", (0 + 4404) => x"00", (0 + 4405) => x"00", (0 + 4406) => x"00", (0 + 4407) => x"00", (0 + 4408) => x"00", (0 + 4409) => x"00", (0 + 4410) => x"00", (0 + 4411) => x"00", (0 + 4412) => x"00", (0 + 4413) => x"00", (0 + 4414) => x"00", (0 + 4415) => x"00", (0 + 4416) => x"00", (0 + 4417) => x"00", (0 + 4418) => x"00", (0 + 4419) => x"00", (0 + 4420) => x"00", (0 + 4421) => x"00", (0 + 4422) => x"00", (0 + 4423) => x"00", (0 + 4424) => x"00", (0 + 4425) => x"00", (0 + 4426) => x"00", (0 + 4427) => x"00", (0 + 4428) => x"00", (0 + 4429) => x"00", (0 + 4430) => x"00", (0 + 4431) => x"00", (0 + 4432) => x"00", (0 + 4433) => x"00", (0 + 4434) => x"00", (0 + 4435) => x"00", (0 + 4436) => x"00", (0 + 4437) => x"00", (0 + 4438) => x"00", (0 + 4439) => x"00", (0 + 4440) => x"00", (0 + 4441) => x"00", (0 + 4442) => x"00", (0 + 4443) => x"00", (0 + 4444) => x"00", (0 + 4445) => x"00", (0 + 4446) => x"00", (0 + 4447) => x"00", (0 + 4448) => x"00", (0 + 4449) => x"00", (0 + 4450) => x"00", (0 + 4451) => x"00", (0 + 4452) => x"00", (0 + 4453) => x"00", (0 + 4454) => x"00", (0 + 4455) => x"00", (0 + 4456) => x"00", (0 + 4457) => x"00", (0 + 4458) => x"00", (0 + 4459) => x"00", (0 + 4460) => x"00", (0 + 4461) => x"00", (0 + 4462) => x"00", (0 + 4463) => x"00", (0 + 4464) => x"00", (0 + 4465) => x"00", (0 + 4466) => x"00", (0 + 4467) => x"00", (0 + 4468) => x"00", (0 + 4469) => x"00", (0 + 4470) => x"00", (0 + 4471) => x"00", (0 + 4472) => x"00", (0 + 4473) => x"00", (0 + 4474) => x"00", (0 + 4475) => x"00", (0 + 4476) => x"00", (0 + 4477) => x"00", (0 + 4478) => x"00", (0 + 4479) => x"00", (0 + 4480) => x"00", (0 + 4481) => x"00", (0 + 4482) => x"00", (0 + 4483) => x"00", (0 + 4484) => x"00", (0 + 4485) => x"00", (0 + 4486) => x"00", (0 + 4487) => x"00", (0 + 4488) => x"00", (0 + 4489) => x"00", (0 + 4490) => x"00", (0 + 4491) => x"00", (0 + 4492) => x"00", (0 + 4493) => x"00", (0 + 4494) => x"00", (0 + 4495) => x"00", (0 + 4496) => x"00", (0 + 4497) => x"00", (0 + 4498) => x"00", (0 + 4499) => x"00", (0 + 4500) => x"00", (0 + 4501) => x"00", (0 + 4502) => x"00", (0 + 4503) => x"00", (0 + 4504) => x"00", (0 + 4505) => x"00", (0 + 4506) => x"00", (0 + 4507) => x"00", (0 + 4508) => x"00", (0 + 4509) => x"00", (0 + 4510) => x"00", (0 + 4511) => x"00", (0 + 4512) => x"00", (0 + 4513) => x"00", (0 + 4514) => x"00", (0 + 4515) => x"00", (0 + 4516) => x"00", (0 + 4517) => x"00", (0 + 4518) => x"00", (0 + 4519) => x"00", (0 + 4520) => x"00", (0 + 4521) => x"00", (0 + 4522) => x"00", (0 + 4523) => x"00", (0 + 4524) => x"00", (0 + 4525) => x"00", (0 + 4526) => x"00", (0 + 4527) => x"00", (0 + 4528) => x"00", (0 + 4529) => x"00", (0 + 4530) => x"00", (0 + 4531) => x"00", (0 + 4532) => x"00", (0 + 4533) => x"00", (0 + 4534) => x"00", (0 + 4535) => x"00", (0 + 4536) => x"00", (0 + 4537) => x"00", (0 + 4538) => x"00", (0 + 4539) => x"00", (0 + 4540) => x"00", (0 + 4541) => x"00", (0 + 4542) => x"00", (0 + 4543) => x"00", (0 + 4544) => x"00", (0 + 4545) => x"00", (0 + 4546) => x"00", (0 + 4547) => x"00", (0 + 4548) => x"00", (0 + 4549) => x"00", (0 + 4550) => x"00", (0 + 4551) => x"00", (0 + 4552) => x"00", (0 + 4553) => x"00", (0 + 4554) => x"00", (0 + 4555) => x"00", (0 + 4556) => x"00", (0 + 4557) => x"00", (0 + 4558) => x"00", (0 + 4559) => x"00", (0 + 4560) => x"00", (0 + 4561) => x"00", (0 + 4562) => x"00", (0 + 4563) => x"00", (0 + 4564) => x"00", (0 + 4565) => x"00", (0 + 4566) => x"00", (0 + 4567) => x"00", (0 + 4568) => x"00", (0 + 4569) => x"00", (0 + 4570) => x"00", (0 + 4571) => x"00", (0 + 4572) => x"00", (0 + 4573) => x"00", (0 + 4574) => x"00", (0 + 4575) => x"00", (0 + 4576) => x"00", (0 + 4577) => x"00", (0 + 4578) => x"00", (0 + 4579) => x"00", (0 + 4580) => x"00", (0 + 4581) => x"00", (0 + 4582) => x"00", (0 + 4583) => x"00", (0 + 4584) => x"00", (0 + 4585) => x"00", (0 + 4586) => x"00", (0 + 4587) => x"00", (0 + 4588) => x"00", (0 + 4589) => x"00", (0 + 4590) => x"00", (0 + 4591) => x"00", (0 + 4592) => x"00", (0 + 4593) => x"00", (0 + 4594) => x"00", (0 + 4595) => x"00", (0 + 4596) => x"00", (0 + 4597) => x"00", (0 + 4598) => x"00", (0 + 4599) => x"00", (0 + 4600) => x"00", (0 + 4601) => x"00", (0 + 4602) => x"00", (0 + 4603) => x"00", (0 + 4604) => x"00", (0 + 4605) => x"00", (0 + 4606) => x"00", (0 + 4607) => x"00", (0 + 4608) => x"00", (0 + 4609) => x"00", (0 + 4610) => x"00", (0 + 4611) => x"00", (0 + 4612) => x"00", (0 + 4613) => x"00", (0 + 4614) => x"00", (0 + 4615) => x"00", (0 + 4616) => x"00", (0 + 4617) => x"00", (0 + 4618) => x"00", (0 + 4619) => x"00", (0 + 4620) => x"00", (0 + 4621) => x"00", (0 + 4622) => x"00", (0 + 4623) => x"00", (0 + 4624) => x"00", (0 + 4625) => x"00", (0 + 4626) => x"00", (0 + 4627) => x"00", (0 + 4628) => x"00", (0 + 4629) => x"00", (0 + 4630) => x"00", (0 + 4631) => x"00", (0 + 4632) => x"00", (0 + 4633) => x"00", (0 + 4634) => x"00", (0 + 4635) => x"00", (0 + 4636) => x"00", (0 + 4637) => x"00", (0 + 4638) => x"00", (0 + 4639) => x"00", (0 + 4640) => x"00", (0 + 4641) => x"00", (0 + 4642) => x"00", (0 + 4643) => x"00", (0 + 4644) => x"00", (0 + 4645) => x"00", (0 + 4646) => x"00", (0 + 4647) => x"00", (0 + 4648) => x"00", (0 + 4649) => x"00", (0 + 4650) => x"00", (0 + 4651) => x"00", (0 + 4652) => x"00", (0 + 4653) => x"00", (0 + 4654) => x"00", (0 + 4655) => x"00", (0 + 4656) => x"00", (0 + 4657) => x"00", (0 + 4658) => x"00", (0 + 4659) => x"00", (0 + 4660) => x"00", (0 + 4661) => x"00", (0 + 4662) => x"00", (0 + 4663) => x"00", (0 + 4664) => x"00", (0 + 4665) => x"00", (0 + 4666) => x"00", (0 + 4667) => x"00", (0 + 4668) => x"00", (0 + 4669) => x"00", (0 + 4670) => x"00", (0 + 4671) => x"00", (0 + 4672) => x"00", (0 + 4673) => x"00", (0 + 4674) => x"00", (0 + 4675) => x"00", (0 + 4676) => x"00", (0 + 4677) => x"00", (0 + 4678) => x"00", (0 + 4679) => x"00", (0 + 4680) => x"00", (0 + 4681) => x"00", (0 + 4682) => x"00", (0 + 4683) => x"00", (0 + 4684) => x"00", (0 + 4685) => x"00", (0 + 4686) => x"00", (0 + 4687) => x"00", (0 + 4688) => x"00", (0 + 4689) => x"00", (0 + 4690) => x"00", (0 + 4691) => x"00", (0 + 4692) => x"00", (0 + 4693) => x"00", (0 + 4694) => x"00", (0 + 4695) => x"00", (0 + 4696) => x"00", (0 + 4697) => x"00", (0 + 4698) => x"00", (0 + 4699) => x"00", (0 + 4700) => x"00", (0 + 4701) => x"00", (0 + 4702) => x"00", (0 + 4703) => x"00", (0 + 4704) => x"00", (0 + 4705) => x"00", (0 + 4706) => x"00", (0 + 4707) => x"00", (0 + 4708) => x"00", (0 + 4709) => x"00", (0 + 4710) => x"00", (0 + 4711) => x"00", (0 + 4712) => x"00", (0 + 4713) => x"00", (0 + 4714) => x"00", (0 + 4715) => x"00", (0 + 4716) => x"00", (0 + 4717) => x"00", (0 + 4718) => x"00", (0 + 4719) => x"00", (0 + 4720) => x"00", (0 + 4721) => x"00", (0 + 4722) => x"00", (0 + 4723) => x"00", (0 + 4724) => x"00", (0 + 4725) => x"00", (0 + 4726) => x"00", (0 + 4727) => x"00", (0 + 4728) => x"00", (0 + 4729) => x"00", (0 + 4730) => x"00", (0 + 4731) => x"00", (0 + 4732) => x"00", (0 + 4733) => x"00", (0 + 4734) => x"00", (0 + 4735) => x"00", (0 + 4736) => x"00", (0 + 4737) => x"00", (0 + 4738) => x"00", (0 + 4739) => x"00", (0 + 4740) => x"00", (0 + 4741) => x"00", (0 + 4742) => x"00", (0 + 4743) => x"00", (0 + 4744) => x"00", (0 + 4745) => x"00", (0 + 4746) => x"00", (0 + 4747) => x"00", (0 + 4748) => x"00", (0 + 4749) => x"00", (0 + 4750) => x"00", (0 + 4751) => x"00", (0 + 4752) => x"00", (0 + 4753) => x"00", (0 + 4754) => x"00", (0 + 4755) => x"00", (0 + 4756) => x"00", (0 + 4757) => x"00", (0 + 4758) => x"00", (0 + 4759) => x"00", (0 + 4760) => x"00", (0 + 4761) => x"00", (0 + 4762) => x"00", (0 + 4763) => x"00", (0 + 4764) => x"00", (0 + 4765) => x"00", (0 + 4766) => x"00", (0 + 4767) => x"00", (0 + 4768) => x"00", (0 + 4769) => x"00", (0 + 4770) => x"00", (0 + 4771) => x"00", (0 + 4772) => x"00", (0 + 4773) => x"00", (0 + 4774) => x"00", (0 + 4775) => x"00", (0 + 4776) => x"00", (0 + 4777) => x"00", (0 + 4778) => x"00", (0 + 4779) => x"00", (0 + 4780) => x"00", (0 + 4781) => x"00", (0 + 4782) => x"00", (0 + 4783) => x"00", (0 + 4784) => x"00", (0 + 4785) => x"00", (0 + 4786) => x"00", (0 + 4787) => x"00", (0 + 4788) => x"00", (0 + 4789) => x"00", (0 + 4790) => x"00", (0 + 4791) => x"00", (0 + 4792) => x"00", (0 + 4793) => x"00", (0 + 4794) => x"00", (0 + 4795) => x"00", (0 + 4796) => x"00", (0 + 4797) => x"00", (0 + 4798) => x"00", (0 + 4799) => x"00", (0 + 4800) => x"00", (0 + 4801) => x"00", (0 + 4802) => x"00", (0 + 4803) => x"00", (0 + 4804) => x"00", (0 + 4805) => x"00", (0 + 4806) => x"00", (0 + 4807) => x"00", (0 + 4808) => x"00", (0 + 4809) => x"00", (0 + 4810) => x"00", (0 + 4811) => x"00", (0 + 4812) => x"00", (0 + 4813) => x"00", (0 + 4814) => x"00", (0 + 4815) => x"00", (0 + 4816) => x"00", (0 + 4817) => x"00", (0 + 4818) => x"00", (0 + 4819) => x"00", (0 + 4820) => x"00", (0 + 4821) => x"00", (0 + 4822) => x"00", (0 + 4823) => x"00", (0 + 4824) => x"00", (0 + 4825) => x"00", (0 + 4826) => x"00", (0 + 4827) => x"00", (0 + 4828) => x"00", (0 + 4829) => x"00", (0 + 4830) => x"00", (0 + 4831) => x"00", (0 + 4832) => x"00", (0 + 4833) => x"00", (0 + 4834) => x"00", (0 + 4835) => x"00", (0 + 4836) => x"00", (0 + 4837) => x"00", (0 + 4838) => x"00", (0 + 4839) => x"00", (0 + 4840) => x"00", (0 + 4841) => x"00", (0 + 4842) => x"00", (0 + 4843) => x"00", (0 + 4844) => x"00", (0 + 4845) => x"00", (0 + 4846) => x"00", (0 + 4847) => x"00", (0 + 4848) => x"00", (0 + 4849) => x"00", (0 + 4850) => x"00", (0 + 4851) => x"00", (0 + 4852) => x"00", (0 + 4853) => x"00", (0 + 4854) => x"00", (0 + 4855) => x"00", (0 + 4856) => x"00", (0 + 4857) => x"00", (0 + 4858) => x"00", (0 + 4859) => x"00", (0 + 4860) => x"00", (0 + 4861) => x"00", (0 + 4862) => x"00", (0 + 4863) => x"00", (0 + 4864) => x"00", (0 + 4865) => x"00", (0 + 4866) => x"00", (0 + 4867) => x"00", (0 + 4868) => x"00", (0 + 4869) => x"00", (0 + 4870) => x"00", (0 + 4871) => x"00", (0 + 4872) => x"00", (0 + 4873) => x"00", (0 + 4874) => x"00", (0 + 4875) => x"00", (0 + 4876) => x"00", (0 + 4877) => x"00", (0 + 4878) => x"00", (0 + 4879) => x"00", (0 + 4880) => x"00", (0 + 4881) => x"00", (0 + 4882) => x"00", (0 + 4883) => x"00", (0 + 4884) => x"00", (0 + 4885) => x"00", (0 + 4886) => x"00", (0 + 4887) => x"00", (0 + 4888) => x"00", (0 + 4889) => x"00", (0 + 4890) => x"00", (0 + 4891) => x"00", (0 + 4892) => x"00", (0 + 4893) => x"00", (0 + 4894) => x"00", (0 + 4895) => x"00", (0 + 4896) => x"00", (0 + 4897) => x"00", (0 + 4898) => x"00", (0 + 4899) => x"00", (0 + 4900) => x"00", (0 + 4901) => x"00", (0 + 4902) => x"00", (0 + 4903) => x"00", (0 + 4904) => x"00", (0 + 4905) => x"00", (0 + 4906) => x"00", (0 + 4907) => x"00", (0 + 4908) => x"00", (0 + 4909) => x"00", (0 + 4910) => x"00", (0 + 4911) => x"00", (0 + 4912) => x"00", (0 + 4913) => x"00", (0 + 4914) => x"00", (0 + 4915) => x"00", (0 + 4916) => x"00", (0 + 4917) => x"00", (0 + 4918) => x"00", (0 + 4919) => x"00", (0 + 4920) => x"00", (0 + 4921) => x"00", (0 + 4922) => x"00", (0 + 4923) => x"00", (0 + 4924) => x"00", (0 + 4925) => x"00", (0 + 4926) => x"00", (0 + 4927) => x"00", (0 + 4928) => x"00", (0 + 4929) => x"00", (0 + 4930) => x"00", (0 + 4931) => x"00", (0 + 4932) => x"00", (0 + 4933) => x"00", (0 + 4934) => x"00", (0 + 4935) => x"00", (0 + 4936) => x"00", (0 + 4937) => x"00", (0 + 4938) => x"00", (0 + 4939) => x"00", (0 + 4940) => x"00", (0 + 4941) => x"00", (0 + 4942) => x"00", (0 + 4943) => x"00", (0 + 4944) => x"00", (0 + 4945) => x"00", (0 + 4946) => x"00", (0 + 4947) => x"00", (0 + 4948) => x"00", (0 + 4949) => x"00", (0 + 4950) => x"00", (0 + 4951) => x"00", (0 + 4952) => x"00", (0 + 4953) => x"00", (0 + 4954) => x"00", (0 + 4955) => x"00", (0 + 4956) => x"00", (0 + 4957) => x"00", (0 + 4958) => x"00", (0 + 4959) => x"00", (0 + 4960) => x"00", (0 + 4961) => x"00", (0 + 4962) => x"00", (0 + 4963) => x"00", (0 + 4964) => x"00", (0 + 4965) => x"00", (0 + 4966) => x"00", (0 + 4967) => x"00", (0 + 4968) => x"00", (0 + 4969) => x"00", (0 + 4970) => x"00", (0 + 4971) => x"00", (0 + 4972) => x"00", (0 + 4973) => x"00", (0 + 4974) => x"00", (0 + 4975) => x"00", (0 + 4976) => x"00", (0 + 4977) => x"00", (0 + 4978) => x"00", (0 + 4979) => x"00", (0 + 4980) => x"00", (0 + 4981) => x"00", (0 + 4982) => x"00", (0 + 4983) => x"00", (0 + 4984) => x"00", (0 + 4985) => x"00", (0 + 4986) => x"00", (0 + 4987) => x"00", (0 + 4988) => x"00", (0 + 4989) => x"00", (0 + 4990) => x"00", (0 + 4991) => x"00", (0 + 4992) => x"00", (0 + 4993) => x"00", (0 + 4994) => x"00", (0 + 4995) => x"00", (0 + 4996) => x"00", (0 + 4997) => x"00", (0 + 4998) => x"00", (0 + 4999) => x"00", (0 + 5000) => x"00", (0 + 5001) => x"00", (0 + 5002) => x"00", (0 + 5003) => x"00", (0 + 5004) => x"00", (0 + 5005) => x"00", (0 + 5006) => x"00", (0 + 5007) => x"00", (0 + 5008) => x"00", (0 + 5009) => x"00", (0 + 5010) => x"00", (0 + 5011) => x"00", (0 + 5012) => x"00", (0 + 5013) => x"00", (0 + 5014) => x"00", (0 + 5015) => x"00", (0 + 5016) => x"00", (0 + 5017) => x"00", (0 + 5018) => x"00", (0 + 5019) => x"00", (0 + 5020) => x"00", (0 + 5021) => x"00", (0 + 5022) => x"00", (0 + 5023) => x"00", (0 + 5024) => x"00", (0 + 5025) => x"00", (0 + 5026) => x"00", (0 + 5027) => x"00", (0 + 5028) => x"00", (0 + 5029) => x"00", (0 + 5030) => x"00", (0 + 5031) => x"00", (0 + 5032) => x"00", (0 + 5033) => x"00", (0 + 5034) => x"00", (0 + 5035) => x"00", (0 + 5036) => x"00", (0 + 5037) => x"00", (0 + 5038) => x"00", (0 + 5039) => x"00", (0 + 5040) => x"00", (0 + 5041) => x"00", (0 + 5042) => x"00", (0 + 5043) => x"00", (0 + 5044) => x"00", (0 + 5045) => x"00", (0 + 5046) => x"00", (0 + 5047) => x"00", (0 + 5048) => x"00", (0 + 5049) => x"00", (0 + 5050) => x"00", (0 + 5051) => x"00", (0 + 5052) => x"00", (0 + 5053) => x"00", (0 + 5054) => x"00", (0 + 5055) => x"00", (0 + 5056) => x"00", (0 + 5057) => x"00", (0 + 5058) => x"00", (0 + 5059) => x"00", (0 + 5060) => x"00", (0 + 5061) => x"00", (0 + 5062) => x"00", (0 + 5063) => x"00", (0 + 5064) => x"00", (0 + 5065) => x"00", (0 + 5066) => x"00", (0 + 5067) => x"00", (0 + 5068) => x"00", (0 + 5069) => x"00", (0 + 5070) => x"00", (0 + 5071) => x"00", (0 + 5072) => x"00", (0 + 5073) => x"00", (0 + 5074) => x"00", (0 + 5075) => x"00", (0 + 5076) => x"00", (0 + 5077) => x"00", (0 + 5078) => x"00", (0 + 5079) => x"00", (0 + 5080) => x"00", (0 + 5081) => x"00", (0 + 5082) => x"00", (0 + 5083) => x"00", (0 + 5084) => x"00", (0 + 5085) => x"00", (0 + 5086) => x"00", (0 + 5087) => x"00", (0 + 5088) => x"00", (0 + 5089) => x"00", (0 + 5090) => x"00", (0 + 5091) => x"00", (0 + 5092) => x"00", (0 + 5093) => x"00", (0 + 5094) => x"00", (0 + 5095) => x"00", (0 + 5096) => x"00", (0 + 5097) => x"00", (0 + 5098) => x"00", (0 + 5099) => x"00", (0 + 5100) => x"00", (0 + 5101) => x"00", (0 + 5102) => x"00", (0 + 5103) => x"00", (0 + 5104) => x"00", (0 + 5105) => x"00", (0 + 5106) => x"00", (0 + 5107) => x"00", (0 + 5108) => x"00", (0 + 5109) => x"00", (0 + 5110) => x"00", (0 + 5111) => x"00", (0 + 5112) => x"00", (0 + 5113) => x"00", (0 + 5114) => x"00", (0 + 5115) => x"00", (0 + 5116) => x"00", (0 + 5117) => x"00", (0 + 5118) => x"00", (0 + 5119) => x"00", (0 + 5120) => x"00", (0 + 5121) => x"00", (0 + 5122) => x"00", (0 + 5123) => x"00", (0 + 5124) => x"00", (0 + 5125) => x"00", (0 + 5126) => x"00", (0 + 5127) => x"00", (0 + 5128) => x"00", (0 + 5129) => x"00", (0 + 5130) => x"00", (0 + 5131) => x"00", (0 + 5132) => x"00", (0 + 5133) => x"00", (0 + 5134) => x"00", (0 + 5135) => x"00", (0 + 5136) => x"00", (0 + 5137) => x"00", (0 + 5138) => x"00", (0 + 5139) => x"00", (0 + 5140) => x"00", (0 + 5141) => x"00", (0 + 5142) => x"00", (0 + 5143) => x"00", (0 + 5144) => x"00", (0 + 5145) => x"00", (0 + 5146) => x"00", (0 + 5147) => x"00", (0 + 5148) => x"00", (0 + 5149) => x"00", (0 + 5150) => x"00", (0 + 5151) => x"00", (0 + 5152) => x"00", (0 + 5153) => x"00", (0 + 5154) => x"00", (0 + 5155) => x"00", (0 + 5156) => x"00", (0 + 5157) => x"00", (0 + 5158) => x"00", (0 + 5159) => x"00", (0 + 5160) => x"00", (0 + 5161) => x"00", (0 + 5162) => x"00", (0 + 5163) => x"00", (0 + 5164) => x"00", (0 + 5165) => x"00", (0 + 5166) => x"00", (0 + 5167) => x"00", (0 + 5168) => x"00", (0 + 5169) => x"00", (0 + 5170) => x"00", (0 + 5171) => x"00", (0 + 5172) => x"00", (0 + 5173) => x"00", (0 + 5174) => x"00", (0 + 5175) => x"00", (0 + 5176) => x"00", (0 + 5177) => x"00", (0 + 5178) => x"00", (0 + 5179) => x"00", (0 + 5180) => x"00", (0 + 5181) => x"00", (0 + 5182) => x"00", (0 + 5183) => x"00", (0 + 5184) => x"00", (0 + 5185) => x"00", (0 + 5186) => x"00", (0 + 5187) => x"00", (0 + 5188) => x"00", (0 + 5189) => x"00", (0 + 5190) => x"00", (0 + 5191) => x"00", (0 + 5192) => x"00", (0 + 5193) => x"00", (0 + 5194) => x"00", (0 + 5195) => x"00", (0 + 5196) => x"00", (0 + 5197) => x"00", (0 + 5198) => x"00", (0 + 5199) => x"00", (0 + 5200) => x"00", (0 + 5201) => x"00", (0 + 5202) => x"00", (0 + 5203) => x"00", (0 + 5204) => x"00", (0 + 5205) => x"00", (0 + 5206) => x"00", (0 + 5207) => x"00", (0 + 5208) => x"00", (0 + 5209) => x"00", (0 + 5210) => x"00", (0 + 5211) => x"00", (0 + 5212) => x"00", (0 + 5213) => x"00", (0 + 5214) => x"00", (0 + 5215) => x"00", (0 + 5216) => x"00", (0 + 5217) => x"00", (0 + 5218) => x"00", (0 + 5219) => x"00", (0 + 5220) => x"00", (0 + 5221) => x"00", (0 + 5222) => x"00", (0 + 5223) => x"00", (0 + 5224) => x"00", (0 + 5225) => x"00", (0 + 5226) => x"00", (0 + 5227) => x"00", (0 + 5228) => x"00", (0 + 5229) => x"00", (0 + 5230) => x"00", (0 + 5231) => x"00", (0 + 5232) => x"00", (0 + 5233) => x"00", (0 + 5234) => x"00", (0 + 5235) => x"00", (0 + 5236) => x"00", (0 + 5237) => x"00", (0 + 5238) => x"00", (0 + 5239) => x"00", (0 + 5240) => x"00", (0 + 5241) => x"00", (0 + 5242) => x"00", (0 + 5243) => x"00", (0 + 5244) => x"00", (0 + 5245) => x"00", (0 + 5246) => x"00", (0 + 5247) => x"00", (0 + 5248) => x"00", (0 + 5249) => x"00", (0 + 5250) => x"00", (0 + 5251) => x"00", (0 + 5252) => x"00", (0 + 5253) => x"00", (0 + 5254) => x"00", (0 + 5255) => x"00", (0 + 5256) => x"00", (0 + 5257) => x"00", (0 + 5258) => x"00", (0 + 5259) => x"00", (0 + 5260) => x"00", (0 + 5261) => x"00", (0 + 5262) => x"00", (0 + 5263) => x"00", (0 + 5264) => x"00", (0 + 5265) => x"00", (0 + 5266) => x"00", (0 + 5267) => x"00", (0 + 5268) => x"00", (0 + 5269) => x"00", (0 + 5270) => x"00", (0 + 5271) => x"00", (0 + 5272) => x"00", (0 + 5273) => x"00", (0 + 5274) => x"00", (0 + 5275) => x"00", (0 + 5276) => x"00", (0 + 5277) => x"00", (0 + 5278) => x"00", (0 + 5279) => x"00", (0 + 5280) => x"00", (0 + 5281) => x"00", (0 + 5282) => x"00", (0 + 5283) => x"00", (0 + 5284) => x"00", (0 + 5285) => x"00", (0 + 5286) => x"00", (0 + 5287) => x"00", (0 + 5288) => x"00", (0 + 5289) => x"00", (0 + 5290) => x"00", (0 + 5291) => x"00", (0 + 5292) => x"00", (0 + 5293) => x"00", (0 + 5294) => x"00", (0 + 5295) => x"00", (0 + 5296) => x"00", (0 + 5297) => x"00", (0 + 5298) => x"00", (0 + 5299) => x"00", (0 + 5300) => x"00", (0 + 5301) => x"00", (0 + 5302) => x"00", (0 + 5303) => x"00", (0 + 5304) => x"00", (0 + 5305) => x"00", (0 + 5306) => x"00", (0 + 5307) => x"00", (0 + 5308) => x"00", (0 + 5309) => x"00", (0 + 5310) => x"00", (0 + 5311) => x"00", (0 + 5312) => x"00", (0 + 5313) => x"00", (0 + 5314) => x"00", (0 + 5315) => x"00", (0 + 5316) => x"00", (0 + 5317) => x"00", (0 + 5318) => x"00", (0 + 5319) => x"00", (0 + 5320) => x"00", (0 + 5321) => x"00", (0 + 5322) => x"00", (0 + 5323) => x"00", (0 + 5324) => x"00", (0 + 5325) => x"00", (0 + 5326) => x"00", (0 + 5327) => x"00", (0 + 5328) => x"00", (0 + 5329) => x"00", (0 + 5330) => x"00", (0 + 5331) => x"00", (0 + 5332) => x"00", (0 + 5333) => x"00", (0 + 5334) => x"00", (0 + 5335) => x"00", (0 + 5336) => x"00", (0 + 5337) => x"00", (0 + 5338) => x"00", (0 + 5339) => x"00", (0 + 5340) => x"00", (0 + 5341) => x"00", (0 + 5342) => x"00", (0 + 5343) => x"00", (0 + 5344) => x"00", (0 + 5345) => x"00", (0 + 5346) => x"00", (0 + 5347) => x"00", (0 + 5348) => x"00", (0 + 5349) => x"00", (0 + 5350) => x"00", (0 + 5351) => x"00", (0 + 5352) => x"00", (0 + 5353) => x"00", (0 + 5354) => x"00", (0 + 5355) => x"00", (0 + 5356) => x"00", (0 + 5357) => x"00", (0 + 5358) => x"00", (0 + 5359) => x"00", (0 + 5360) => x"00", (0 + 5361) => x"00", (0 + 5362) => x"00", (0 + 5363) => x"00", (0 + 5364) => x"00", (0 + 5365) => x"00", (0 + 5366) => x"00", (0 + 5367) => x"00", (0 + 5368) => x"00", (0 + 5369) => x"00", (0 + 5370) => x"00", (0 + 5371) => x"00", (0 + 5372) => x"00", (0 + 5373) => x"00", (0 + 5374) => x"00", (0 + 5375) => x"00", (0 + 5376) => x"00", (0 + 5377) => x"00", (0 + 5378) => x"00", (0 + 5379) => x"00", (0 + 5380) => x"00", (0 + 5381) => x"00", (0 + 5382) => x"00", (0 + 5383) => x"00", (0 + 5384) => x"00", (0 + 5385) => x"00", (0 + 5386) => x"00", (0 + 5387) => x"00", (0 + 5388) => x"00", (0 + 5389) => x"00", (0 + 5390) => x"00", (0 + 5391) => x"00", (0 + 5392) => x"00", (0 + 5393) => x"00", (0 + 5394) => x"00", (0 + 5395) => x"00", (0 + 5396) => x"00", (0 + 5397) => x"00", (0 + 5398) => x"00", (0 + 5399) => x"00", (0 + 5400) => x"00", (0 + 5401) => x"00", (0 + 5402) => x"00", (0 + 5403) => x"00", (0 + 5404) => x"00", (0 + 5405) => x"00", (0 + 5406) => x"00", (0 + 5407) => x"00", (0 + 5408) => x"00", (0 + 5409) => x"00", (0 + 5410) => x"00", (0 + 5411) => x"00", (0 + 5412) => x"00", (0 + 5413) => x"00", (0 + 5414) => x"00", (0 + 5415) => x"00", (0 + 5416) => x"00", (0 + 5417) => x"00", (0 + 5418) => x"00", (0 + 5419) => x"00", (0 + 5420) => x"00", (0 + 5421) => x"00", (0 + 5422) => x"00", (0 + 5423) => x"00", (0 + 5424) => x"00", (0 + 5425) => x"00", (0 + 5426) => x"00", (0 + 5427) => x"00", (0 + 5428) => x"00", (0 + 5429) => x"00", (0 + 5430) => x"00", (0 + 5431) => x"00", (0 + 5432) => x"00", (0 + 5433) => x"00", (0 + 5434) => x"00", (0 + 5435) => x"00", (0 + 5436) => x"00", (0 + 5437) => x"00", (0 + 5438) => x"00", (0 + 5439) => x"00", (0 + 5440) => x"00", (0 + 5441) => x"00", (0 + 5442) => x"00", (0 + 5443) => x"00", (0 + 5444) => x"00", (0 + 5445) => x"00", (0 + 5446) => x"00", (0 + 5447) => x"00", (0 + 5448) => x"00", (0 + 5449) => x"00", (0 + 5450) => x"00", (0 + 5451) => x"00", (0 + 5452) => x"00", (0 + 5453) => x"00", (0 + 5454) => x"00", (0 + 5455) => x"00", (0 + 5456) => x"00", (0 + 5457) => x"00", (0 + 5458) => x"00", (0 + 5459) => x"00", (0 + 5460) => x"00", (0 + 5461) => x"00", (0 + 5462) => x"00", (0 + 5463) => x"00", (0 + 5464) => x"00", (0 + 5465) => x"00", (0 + 5466) => x"00", (0 + 5467) => x"00", (0 + 5468) => x"00", (0 + 5469) => x"00", (0 + 5470) => x"00", (0 + 5471) => x"00", (0 + 5472) => x"00", (0 + 5473) => x"00", (0 + 5474) => x"00", (0 + 5475) => x"00", (0 + 5476) => x"00", (0 + 5477) => x"00", (0 + 5478) => x"00", (0 + 5479) => x"00", (0 + 5480) => x"00", (0 + 5481) => x"00", (0 + 5482) => x"00", (0 + 5483) => x"00", (0 + 5484) => x"00", (0 + 5485) => x"00", (0 + 5486) => x"00", (0 + 5487) => x"00", (0 + 5488) => x"00", (0 + 5489) => x"00", (0 + 5490) => x"00", (0 + 5491) => x"00", (0 + 5492) => x"00", (0 + 5493) => x"00", (0 + 5494) => x"00", (0 + 5495) => x"00", (0 + 5496) => x"00", (0 + 5497) => x"00", (0 + 5498) => x"00", (0 + 5499) => x"00", (0 + 5500) => x"00", (0 + 5501) => x"00", (0 + 5502) => x"00", (0 + 5503) => x"00", (0 + 5504) => x"00", (0 + 5505) => x"00", (0 + 5506) => x"00", (0 + 5507) => x"00", (0 + 5508) => x"00", (0 + 5509) => x"00", (0 + 5510) => x"00", (0 + 5511) => x"00", (0 + 5512) => x"00", (0 + 5513) => x"00", (0 + 5514) => x"00", (0 + 5515) => x"00", (0 + 5516) => x"00", (0 + 5517) => x"00", (0 + 5518) => x"00", (0 + 5519) => x"00", (0 + 5520) => x"00", (0 + 5521) => x"00", (0 + 5522) => x"00", (0 + 5523) => x"00", (0 + 5524) => x"00", (0 + 5525) => x"00", (0 + 5526) => x"00", (0 + 5527) => x"00", (0 + 5528) => x"00", (0 + 5529) => x"00", (0 + 5530) => x"00", (0 + 5531) => x"00", (0 + 5532) => x"00", (0 + 5533) => x"00", (0 + 5534) => x"00", (0 + 5535) => x"00", (0 + 5536) => x"00", (0 + 5537) => x"00", (0 + 5538) => x"00", (0 + 5539) => x"00", (0 + 5540) => x"00", (0 + 5541) => x"00", (0 + 5542) => x"00", (0 + 5543) => x"00", (0 + 5544) => x"00", (0 + 5545) => x"00", (0 + 5546) => x"00", (0 + 5547) => x"00", (0 + 5548) => x"00", (0 + 5549) => x"00", (0 + 5550) => x"00", (0 + 5551) => x"00", (0 + 5552) => x"00", (0 + 5553) => x"00", (0 + 5554) => x"00", (0 + 5555) => x"00", (0 + 5556) => x"00", (0 + 5557) => x"00", (0 + 5558) => x"00", (0 + 5559) => x"00", (0 + 5560) => x"00", (0 + 5561) => x"00", (0 + 5562) => x"00", (0 + 5563) => x"00", (0 + 5564) => x"00", (0 + 5565) => x"00", (0 + 5566) => x"00", (0 + 5567) => x"00", (0 + 5568) => x"00", (0 + 5569) => x"00", (0 + 5570) => x"00", (0 + 5571) => x"00", (0 + 5572) => x"00", (0 + 5573) => x"00", (0 + 5574) => x"00", (0 + 5575) => x"00", (0 + 5576) => x"00", (0 + 5577) => x"00", (0 + 5578) => x"00", (0 + 5579) => x"00", (0 + 5580) => x"00", (0 + 5581) => x"00", (0 + 5582) => x"00", (0 + 5583) => x"00", (0 + 5584) => x"00", (0 + 5585) => x"00", (0 + 5586) => x"00", (0 + 5587) => x"00", (0 + 5588) => x"00", (0 + 5589) => x"00", (0 + 5590) => x"00", (0 + 5591) => x"00", (0 + 5592) => x"00", (0 + 5593) => x"00", (0 + 5594) => x"00", (0 + 5595) => x"00", (0 + 5596) => x"00", (0 + 5597) => x"00", (0 + 5598) => x"00", (0 + 5599) => x"00", (0 + 5600) => x"00", (0 + 5601) => x"00", (0 + 5602) => x"00", (0 + 5603) => x"00", (0 + 5604) => x"00", (0 + 5605) => x"00", (0 + 5606) => x"00", (0 + 5607) => x"00", (0 + 5608) => x"00", (0 + 5609) => x"00", (0 + 5610) => x"00", (0 + 5611) => x"00", (0 + 5612) => x"00", (0 + 5613) => x"00", (0 + 5614) => x"00", (0 + 5615) => x"00", (0 + 5616) => x"00", (0 + 5617) => x"00", (0 + 5618) => x"00", (0 + 5619) => x"00", (0 + 5620) => x"00", (0 + 5621) => x"00", (0 + 5622) => x"00", (0 + 5623) => x"00", (0 + 5624) => x"00", (0 + 5625) => x"00", (0 + 5626) => x"00", (0 + 5627) => x"00", (0 + 5628) => x"00", (0 + 5629) => x"00", (0 + 5630) => x"00", (0 + 5631) => x"00", (0 + 5632) => x"00", (0 + 5633) => x"00", (0 + 5634) => x"00", (0 + 5635) => x"00", (0 + 5636) => x"00", (0 + 5637) => x"00", (0 + 5638) => x"00", (0 + 5639) => x"00", (0 + 5640) => x"00", (0 + 5641) => x"00", (0 + 5642) => x"00", (0 + 5643) => x"00", (0 + 5644) => x"00", (0 + 5645) => x"00", (0 + 5646) => x"00", (0 + 5647) => x"00", (0 + 5648) => x"00", (0 + 5649) => x"00", (0 + 5650) => x"00", (0 + 5651) => x"00", (0 + 5652) => x"00", (0 + 5653) => x"00", (0 + 5654) => x"00", (0 + 5655) => x"00", (0 + 5656) => x"00", (0 + 5657) => x"00", (0 + 5658) => x"00", (0 + 5659) => x"00", (0 + 5660) => x"00", (0 + 5661) => x"00", (0 + 5662) => x"00", (0 + 5663) => x"00", (0 + 5664) => x"00", (0 + 5665) => x"00", (0 + 5666) => x"00", (0 + 5667) => x"00", (0 + 5668) => x"00", (0 + 5669) => x"00", (0 + 5670) => x"00", (0 + 5671) => x"00", (0 + 5672) => x"00", (0 + 5673) => x"00", (0 + 5674) => x"00", (0 + 5675) => x"00", (0 + 5676) => x"00", (0 + 5677) => x"00", (0 + 5678) => x"00", (0 + 5679) => x"00", (0 + 5680) => x"00", (0 + 5681) => x"00", (0 + 5682) => x"00", (0 + 5683) => x"00", (0 + 5684) => x"00", (0 + 5685) => x"00", (0 + 5686) => x"00", (0 + 5687) => x"00", (0 + 5688) => x"00", (0 + 5689) => x"00", (0 + 5690) => x"00", (0 + 5691) => x"00", (0 + 5692) => x"00", (0 + 5693) => x"00", (0 + 5694) => x"00", (0 + 5695) => x"00", (0 + 5696) => x"00", (0 + 5697) => x"00", (0 + 5698) => x"00", (0 + 5699) => x"00", (0 + 5700) => x"00", (0 + 5701) => x"00", (0 + 5702) => x"00", (0 + 5703) => x"00", (0 + 5704) => x"00", (0 + 5705) => x"00", (0 + 5706) => x"00", (0 + 5707) => x"00", (0 + 5708) => x"00", (0 + 5709) => x"00", (0 + 5710) => x"00", (0 + 5711) => x"00", (0 + 5712) => x"00", (0 + 5713) => x"00", (0 + 5714) => x"00", (0 + 5715) => x"00", (0 + 5716) => x"00", (0 + 5717) => x"00", (0 + 5718) => x"00", (0 + 5719) => x"00", (0 + 5720) => x"00", (0 + 5721) => x"00", (0 + 5722) => x"00", (0 + 5723) => x"00", (0 + 5724) => x"00", (0 + 5725) => x"00", (0 + 5726) => x"00", (0 + 5727) => x"00", (0 + 5728) => x"00", (0 + 5729) => x"00", (0 + 5730) => x"00", (0 + 5731) => x"00", (0 + 5732) => x"00", (0 + 5733) => x"00", (0 + 5734) => x"00", (0 + 5735) => x"00", (0 + 5736) => x"00", (0 + 5737) => x"00", (0 + 5738) => x"00", (0 + 5739) => x"00", (0 + 5740) => x"00", (0 + 5741) => x"00", (0 + 5742) => x"00", (0 + 5743) => x"00", (0 + 5744) => x"00", (0 + 5745) => x"00", (0 + 5746) => x"00", (0 + 5747) => x"00", (0 + 5748) => x"00", (0 + 5749) => x"00", (0 + 5750) => x"00", (0 + 5751) => x"00", (0 + 5752) => x"00", (0 + 5753) => x"00", (0 + 5754) => x"00", (0 + 5755) => x"00", (0 + 5756) => x"00", (0 + 5757) => x"00", (0 + 5758) => x"00", (0 + 5759) => x"00", (0 + 5760) => x"00", (0 + 5761) => x"00", (0 + 5762) => x"00", (0 + 5763) => x"00", (0 + 5764) => x"00", (0 + 5765) => x"00", (0 + 5766) => x"00", (0 + 5767) => x"00", (0 + 5768) => x"00", (0 + 5769) => x"00", (0 + 5770) => x"00", (0 + 5771) => x"00", (0 + 5772) => x"00", (0 + 5773) => x"00", (0 + 5774) => x"00", (0 + 5775) => x"00", (0 + 5776) => x"00", (0 + 5777) => x"00", (0 + 5778) => x"00", (0 + 5779) => x"00", (0 + 5780) => x"00", (0 + 5781) => x"00", (0 + 5782) => x"00", (0 + 5783) => x"00", (0 + 5784) => x"00", (0 + 5785) => x"00", (0 + 5786) => x"00", (0 + 5787) => x"00", (0 + 5788) => x"00", (0 + 5789) => x"00", (0 + 5790) => x"00", (0 + 5791) => x"00", (0 + 5792) => x"00", (0 + 5793) => x"00", (0 + 5794) => x"00", (0 + 5795) => x"00", (0 + 5796) => x"00", (0 + 5797) => x"00", (0 + 5798) => x"00", (0 + 5799) => x"00", (0 + 5800) => x"00", (0 + 5801) => x"00", (0 + 5802) => x"00", (0 + 5803) => x"00", (0 + 5804) => x"00", (0 + 5805) => x"00", (0 + 5806) => x"00", (0 + 5807) => x"00", (0 + 5808) => x"00", (0 + 5809) => x"00", (0 + 5810) => x"00", (0 + 5811) => x"00", (0 + 5812) => x"00", (0 + 5813) => x"00", (0 + 5814) => x"00", (0 + 5815) => x"00", (0 + 5816) => x"00", (0 + 5817) => x"00", (0 + 5818) => x"00", (0 + 5819) => x"00", (0 + 5820) => x"00", (0 + 5821) => x"00", (0 + 5822) => x"00", (0 + 5823) => x"00", (0 + 5824) => x"00", (0 + 5825) => x"00", (0 + 5826) => x"00", (0 + 5827) => x"00", (0 + 5828) => x"00", (0 + 5829) => x"00", (0 + 5830) => x"00", (0 + 5831) => x"00", (0 + 5832) => x"00", (0 + 5833) => x"00", (0 + 5834) => x"00", (0 + 5835) => x"00", (0 + 5836) => x"00", (0 + 5837) => x"00", (0 + 5838) => x"00", (0 + 5839) => x"00", (0 + 5840) => x"00", (0 + 5841) => x"00", (0 + 5842) => x"00", (0 + 5843) => x"00", (0 + 5844) => x"00", (0 + 5845) => x"00", (0 + 5846) => x"00", (0 + 5847) => x"00", (0 + 5848) => x"00", (0 + 5849) => x"00", (0 + 5850) => x"00", (0 + 5851) => x"00", (0 + 5852) => x"00", (0 + 5853) => x"00", (0 + 5854) => x"00", (0 + 5855) => x"00", (0 + 5856) => x"00", (0 + 5857) => x"00", (0 + 5858) => x"00", (0 + 5859) => x"00", (0 + 5860) => x"00", (0 + 5861) => x"00", (0 + 5862) => x"00", (0 + 5863) => x"00", (0 + 5864) => x"00", (0 + 5865) => x"00", (0 + 5866) => x"00", (0 + 5867) => x"00", (0 + 5868) => x"00", (0 + 5869) => x"00", (0 + 5870) => x"00", (0 + 5871) => x"00", (0 + 5872) => x"00", (0 + 5873) => x"00", (0 + 5874) => x"00", (0 + 5875) => x"00", (0 + 5876) => x"00", (0 + 5877) => x"00", (0 + 5878) => x"00", (0 + 5879) => x"00", (0 + 5880) => x"00", (0 + 5881) => x"00", (0 + 5882) => x"00", (0 + 5883) => x"00", (0 + 5884) => x"00", (0 + 5885) => x"00", (0 + 5886) => x"00", (0 + 5887) => x"00", (0 + 5888) => x"00", (0 + 5889) => x"00", (0 + 5890) => x"00", (0 + 5891) => x"00", (0 + 5892) => x"00", (0 + 5893) => x"00", (0 + 5894) => x"00", (0 + 5895) => x"00", (0 + 5896) => x"00", (0 + 5897) => x"00", (0 + 5898) => x"00", (0 + 5899) => x"00", (0 + 5900) => x"00", (0 + 5901) => x"00", (0 + 5902) => x"00", (0 + 5903) => x"00", (0 + 5904) => x"00", (0 + 5905) => x"00", (0 + 5906) => x"00", (0 + 5907) => x"00", (0 + 5908) => x"00", (0 + 5909) => x"00", (0 + 5910) => x"00", (0 + 5911) => x"00", (0 + 5912) => x"00", (0 + 5913) => x"00", (0 + 5914) => x"00", (0 + 5915) => x"00", (0 + 5916) => x"00", (0 + 5917) => x"00", (0 + 5918) => x"00", (0 + 5919) => x"00", (0 + 5920) => x"00", (0 + 5921) => x"00", (0 + 5922) => x"00", (0 + 5923) => x"00", (0 + 5924) => x"00", (0 + 5925) => x"00", (0 + 5926) => x"00", (0 + 5927) => x"00", (0 + 5928) => x"00", (0 + 5929) => x"00", (0 + 5930) => x"00", (0 + 5931) => x"00", (0 + 5932) => x"00", (0 + 5933) => x"00", (0 + 5934) => x"00", (0 + 5935) => x"00", (0 + 5936) => x"00", (0 + 5937) => x"00", (0 + 5938) => x"00", (0 + 5939) => x"00", (0 + 5940) => x"00", (0 + 5941) => x"00", (0 + 5942) => x"00", (0 + 5943) => x"00", (0 + 5944) => x"00", (0 + 5945) => x"00", (0 + 5946) => x"00", (0 + 5947) => x"00", (0 + 5948) => x"00", (0 + 5949) => x"00", (0 + 5950) => x"00", (0 + 5951) => x"00", (0 + 5952) => x"00", (0 + 5953) => x"00", (0 + 5954) => x"00", (0 + 5955) => x"00", (0 + 5956) => x"00", (0 + 5957) => x"00", (0 + 5958) => x"00", (0 + 5959) => x"00", (0 + 5960) => x"00", (0 + 5961) => x"00", (0 + 5962) => x"00", (0 + 5963) => x"00", (0 + 5964) => x"00", (0 + 5965) => x"00", (0 + 5966) => x"00", (0 + 5967) => x"00", (0 + 5968) => x"00", (0 + 5969) => x"00", (0 + 5970) => x"00", (0 + 5971) => x"00", (0 + 5972) => x"00", (0 + 5973) => x"00", (0 + 5974) => x"00", (0 + 5975) => x"00", (0 + 5976) => x"00", (0 + 5977) => x"00", (0 + 5978) => x"00", (0 + 5979) => x"00", (0 + 5980) => x"00", (0 + 5981) => x"00", (0 + 5982) => x"00", (0 + 5983) => x"00", (0 + 5984) => x"00", (0 + 5985) => x"00", (0 + 5986) => x"00", (0 + 5987) => x"00", (0 + 5988) => x"00", (0 + 5989) => x"00", (0 + 5990) => x"00", (0 + 5991) => x"00", (0 + 5992) => x"00", (0 + 5993) => x"00", (0 + 5994) => x"00", (0 + 5995) => x"00", (0 + 5996) => x"00", (0 + 5997) => x"00", (0 + 5998) => x"00", (0 + 5999) => x"00", (0 + 6000) => x"00", (0 + 6001) => x"00", (0 + 6002) => x"00", (0 + 6003) => x"00", (0 + 6004) => x"00", (0 + 6005) => x"00", (0 + 6006) => x"00", (0 + 6007) => x"00", (0 + 6008) => x"00", (0 + 6009) => x"00", (0 + 6010) => x"00", (0 + 6011) => x"00", (0 + 6012) => x"00", (0 + 6013) => x"00", (0 + 6014) => x"00", (0 + 6015) => x"00", (0 + 6016) => x"00", (0 + 6017) => x"00", (0 + 6018) => x"00", (0 + 6019) => x"00", (0 + 6020) => x"00", (0 + 6021) => x"00", (0 + 6022) => x"00", (0 + 6023) => x"00", (0 + 6024) => x"00", (0 + 6025) => x"00", (0 + 6026) => x"00", (0 + 6027) => x"00", (0 + 6028) => x"00", (0 + 6029) => x"00", (0 + 6030) => x"00", (0 + 6031) => x"00", (0 + 6032) => x"00", (0 + 6033) => x"00", (0 + 6034) => x"00", (0 + 6035) => x"00", (0 + 6036) => x"00", (0 + 6037) => x"00", (0 + 6038) => x"00", (0 + 6039) => x"00", (0 + 6040) => x"00", (0 + 6041) => x"00", (0 + 6042) => x"00", (0 + 6043) => x"00", (0 + 6044) => x"00", (0 + 6045) => x"00", (0 + 6046) => x"00", (0 + 6047) => x"00", (0 + 6048) => x"00", (0 + 6049) => x"00", (0 + 6050) => x"00", (0 + 6051) => x"00", (0 + 6052) => x"00", (0 + 6053) => x"00", (0 + 6054) => x"00", (0 + 6055) => x"00", (0 + 6056) => x"00", (0 + 6057) => x"00", (0 + 6058) => x"00", (0 + 6059) => x"00", (0 + 6060) => x"00", (0 + 6061) => x"00", (0 + 6062) => x"00", (0 + 6063) => x"00", (0 + 6064) => x"00", (0 + 6065) => x"00", (0 + 6066) => x"00", (0 + 6067) => x"00", (0 + 6068) => x"00", (0 + 6069) => x"00", (0 + 6070) => x"00", (0 + 6071) => x"00", (0 + 6072) => x"00", (0 + 6073) => x"00", (0 + 6074) => x"00", (0 + 6075) => x"00", (0 + 6076) => x"00", (0 + 6077) => x"00", (0 + 6078) => x"00", (0 + 6079) => x"00", (0 + 6080) => x"00", (0 + 6081) => x"00", (0 + 6082) => x"00", (0 + 6083) => x"00", (0 + 6084) => x"00", (0 + 6085) => x"00", (0 + 6086) => x"00", (0 + 6087) => x"00", (0 + 6088) => x"00", (0 + 6089) => x"00", (0 + 6090) => x"00", (0 + 6091) => x"00", (0 + 6092) => x"00", (0 + 6093) => x"00", (0 + 6094) => x"00", (0 + 6095) => x"00", (0 + 6096) => x"00", (0 + 6097) => x"00", (0 + 6098) => x"00", (0 + 6099) => x"00", (0 + 6100) => x"00", (0 + 6101) => x"00", (0 + 6102) => x"00", (0 + 6103) => x"00", (0 + 6104) => x"00", (0 + 6105) => x"00", (0 + 6106) => x"00", (0 + 6107) => x"00", (0 + 6108) => x"00", (0 + 6109) => x"00", (0 + 6110) => x"00", (0 + 6111) => x"00", (0 + 6112) => x"00", (0 + 6113) => x"00", (0 + 6114) => x"00", (0 + 6115) => x"00", (0 + 6116) => x"00", (0 + 6117) => x"00", (0 + 6118) => x"00", (0 + 6119) => x"00", (0 + 6120) => x"00", (0 + 6121) => x"00", (0 + 6122) => x"00", (0 + 6123) => x"00", (0 + 6124) => x"00", (0 + 6125) => x"00", (0 + 6126) => x"00", (0 + 6127) => x"00", (0 + 6128) => x"00", (0 + 6129) => x"00", (0 + 6130) => x"00", (0 + 6131) => x"00", (0 + 6132) => x"00", (0 + 6133) => x"00", (0 + 6134) => x"00", (0 + 6135) => x"00", (0 + 6136) => x"00", (0 + 6137) => x"00", (0 + 6138) => x"00", (0 + 6139) => x"00", (0 + 6140) => x"00", (0 + 6141) => x"00", (0 + 6142) => x"00", (0 + 6143) => x"00", (0 + 6144) => x"00", (0 + 6145) => x"00", (0 + 6146) => x"00", (0 + 6147) => x"00", (0 + 6148) => x"00", (0 + 6149) => x"00", (0 + 6150) => x"00", (0 + 6151) => x"00", (0 + 6152) => x"00", (0 + 6153) => x"00", (0 + 6154) => x"00", (0 + 6155) => x"00", (0 + 6156) => x"00", (0 + 6157) => x"00", (0 + 6158) => x"00", (0 + 6159) => x"00", (0 + 6160) => x"00", (0 + 6161) => x"00", (0 + 6162) => x"00", (0 + 6163) => x"00", (0 + 6164) => x"00", (0 + 6165) => x"00", (0 + 6166) => x"00", (0 + 6167) => x"00", (0 + 6168) => x"00", (0 + 6169) => x"00", (0 + 6170) => x"00", (0 + 6171) => x"00", (0 + 6172) => x"00", (0 + 6173) => x"00", (0 + 6174) => x"00", (0 + 6175) => x"00", (0 + 6176) => x"00", (0 + 6177) => x"00", (0 + 6178) => x"00", (0 + 6179) => x"00", (0 + 6180) => x"00", (0 + 6181) => x"00", (0 + 6182) => x"00", (0 + 6183) => x"00", (0 + 6184) => x"00", (0 + 6185) => x"00", (0 + 6186) => x"00", (0 + 6187) => x"00", (0 + 6188) => x"00", (0 + 6189) => x"00", (0 + 6190) => x"00", (0 + 6191) => x"00", (0 + 6192) => x"00", (0 + 6193) => x"00", (0 + 6194) => x"00", (0 + 6195) => x"00", (0 + 6196) => x"00", (0 + 6197) => x"00", (0 + 6198) => x"00", (0 + 6199) => x"00", (0 + 6200) => x"00", (0 + 6201) => x"00", (0 + 6202) => x"00", (0 + 6203) => x"00", (0 + 6204) => x"00", (0 + 6205) => x"00", (0 + 6206) => x"00", (0 + 6207) => x"00", (0 + 6208) => x"00", (0 + 6209) => x"00", (0 + 6210) => x"00", (0 + 6211) => x"00", (0 + 6212) => x"00", (0 + 6213) => x"00", (0 + 6214) => x"00", (0 + 6215) => x"00", (0 + 6216) => x"00", (0 + 6217) => x"00", (0 + 6218) => x"00", (0 + 6219) => x"00", (0 + 6220) => x"00", (0 + 6221) => x"00", (0 + 6222) => x"00", (0 + 6223) => x"00", (0 + 6224) => x"00", (0 + 6225) => x"00", (0 + 6226) => x"00", (0 + 6227) => x"00", (0 + 6228) => x"00", (0 + 6229) => x"00", (0 + 6230) => x"00", (0 + 6231) => x"00", (0 + 6232) => x"00", (0 + 6233) => x"00", (0 + 6234) => x"00", (0 + 6235) => x"00", (0 + 6236) => x"00", (0 + 6237) => x"00", (0 + 6238) => x"00", (0 + 6239) => x"00", (0 + 6240) => x"00", (0 + 6241) => x"00", (0 + 6242) => x"00", (0 + 6243) => x"00", (0 + 6244) => x"00", (0 + 6245) => x"00", (0 + 6246) => x"00", (0 + 6247) => x"00", (0 + 6248) => x"00", (0 + 6249) => x"00", (0 + 6250) => x"00", (0 + 6251) => x"00", (0 + 6252) => x"00", (0 + 6253) => x"00", (0 + 6254) => x"00", (0 + 6255) => x"00", (0 + 6256) => x"00", (0 + 6257) => x"00", (0 + 6258) => x"00", (0 + 6259) => x"00", (0 + 6260) => x"00", (0 + 6261) => x"00", (0 + 6262) => x"00", (0 + 6263) => x"00", (0 + 6264) => x"00", (0 + 6265) => x"00", (0 + 6266) => x"00", (0 + 6267) => x"00", (0 + 6268) => x"00", (0 + 6269) => x"00", (0 + 6270) => x"00", (0 + 6271) => x"00", (0 + 6272) => x"00", (0 + 6273) => x"00", (0 + 6274) => x"00", (0 + 6275) => x"00", (0 + 6276) => x"00", (0 + 6277) => x"00", (0 + 6278) => x"00", (0 + 6279) => x"00", (0 + 6280) => x"00", (0 + 6281) => x"00", (0 + 6282) => x"00", (0 + 6283) => x"00", (0 + 6284) => x"00", (0 + 6285) => x"00", (0 + 6286) => x"00", (0 + 6287) => x"00", (0 + 6288) => x"00", (0 + 6289) => x"00", (0 + 6290) => x"00", (0 + 6291) => x"00", (0 + 6292) => x"00", (0 + 6293) => x"00", (0 + 6294) => x"00", (0 + 6295) => x"00", (0 + 6296) => x"00", (0 + 6297) => x"00", (0 + 6298) => x"00", (0 + 6299) => x"00", (0 + 6300) => x"00", (0 + 6301) => x"00", (0 + 6302) => x"00", (0 + 6303) => x"00", (0 + 6304) => x"00", (0 + 6305) => x"00", (0 + 6306) => x"00", (0 + 6307) => x"00", (0 + 6308) => x"00", (0 + 6309) => x"00", (0 + 6310) => x"00", (0 + 6311) => x"00", (0 + 6312) => x"00", (0 + 6313) => x"00", (0 + 6314) => x"00", (0 + 6315) => x"00", (0 + 6316) => x"00", (0 + 6317) => x"00", (0 + 6318) => x"00", (0 + 6319) => x"00", (0 + 6320) => x"00", (0 + 6321) => x"00", (0 + 6322) => x"00", (0 + 6323) => x"00", (0 + 6324) => x"00", (0 + 6325) => x"00", (0 + 6326) => x"00", (0 + 6327) => x"00", (0 + 6328) => x"00", (0 + 6329) => x"00", (0 + 6330) => x"00", (0 + 6331) => x"00", (0 + 6332) => x"00", (0 + 6333) => x"00", (0 + 6334) => x"00", (0 + 6335) => x"00", (0 + 6336) => x"00", (0 + 6337) => x"00", (0 + 6338) => x"00", (0 + 6339) => x"00", (0 + 6340) => x"00", (0 + 6341) => x"00", (0 + 6342) => x"00", (0 + 6343) => x"00", (0 + 6344) => x"00", (0 + 6345) => x"00", (0 + 6346) => x"00", (0 + 6347) => x"00", (0 + 6348) => x"00", (0 + 6349) => x"00", (0 + 6350) => x"00", (0 + 6351) => x"00", (0 + 6352) => x"00", (0 + 6353) => x"00", (0 + 6354) => x"00", (0 + 6355) => x"00", (0 + 6356) => x"00", (0 + 6357) => x"00", (0 + 6358) => x"00", (0 + 6359) => x"00", (0 + 6360) => x"00", (0 + 6361) => x"00", (0 + 6362) => x"00", (0 + 6363) => x"00", (0 + 6364) => x"00", (0 + 6365) => x"00", (0 + 6366) => x"00", (0 + 6367) => x"00", (0 + 6368) => x"00", (0 + 6369) => x"00", (0 + 6370) => x"00", (0 + 6371) => x"00", (0 + 6372) => x"00", (0 + 6373) => x"00", (0 + 6374) => x"00", (0 + 6375) => x"00", (0 + 6376) => x"00", (0 + 6377) => x"00", (0 + 6378) => x"00", (0 + 6379) => x"00", (0 + 6380) => x"00", (0 + 6381) => x"00", (0 + 6382) => x"00", (0 + 6383) => x"00", (0 + 6384) => x"00", (0 + 6385) => x"00", (0 + 6386) => x"00", (0 + 6387) => x"00", (0 + 6388) => x"00", (0 + 6389) => x"00", (0 + 6390) => x"00", (0 + 6391) => x"00", (0 + 6392) => x"00", (0 + 6393) => x"00", (0 + 6394) => x"00", (0 + 6395) => x"00", (0 + 6396) => x"00", (0 + 6397) => x"00", (0 + 6398) => x"00", (0 + 6399) => x"00", (0 + 6400) => x"00", (0 + 6401) => x"00", (0 + 6402) => x"00", (0 + 6403) => x"00", (0 + 6404) => x"00", (0 + 6405) => x"00", (0 + 6406) => x"00", (0 + 6407) => x"00", (0 + 6408) => x"00", (0 + 6409) => x"00", (0 + 6410) => x"00", (0 + 6411) => x"00", (0 + 6412) => x"00", (0 + 6413) => x"00", (0 + 6414) => x"00", (0 + 6415) => x"00", (0 + 6416) => x"00", (0 + 6417) => x"00", (0 + 6418) => x"00", (0 + 6419) => x"00", (0 + 6420) => x"00", (0 + 6421) => x"00", (0 + 6422) => x"00", (0 + 6423) => x"00", (0 + 6424) => x"00", (0 + 6425) => x"00", (0 + 6426) => x"00", (0 + 6427) => x"00", (0 + 6428) => x"00", (0 + 6429) => x"00", (0 + 6430) => x"00", (0 + 6431) => x"00", (0 + 6432) => x"00", (0 + 6433) => x"00", (0 + 6434) => x"00", (0 + 6435) => x"00", (0 + 6436) => x"00", (0 + 6437) => x"00", (0 + 6438) => x"00", (0 + 6439) => x"00", (0 + 6440) => x"00", (0 + 6441) => x"00", (0 + 6442) => x"00", (0 + 6443) => x"00", (0 + 6444) => x"00", (0 + 6445) => x"00", (0 + 6446) => x"00", (0 + 6447) => x"00", (0 + 6448) => x"00", (0 + 6449) => x"00", (0 + 6450) => x"00", (0 + 6451) => x"00", (0 + 6452) => x"00", (0 + 6453) => x"00", (0 + 6454) => x"00", (0 + 6455) => x"00", (0 + 6456) => x"00", (0 + 6457) => x"00", (0 + 6458) => x"00", (0 + 6459) => x"00", (0 + 6460) => x"00", (0 + 6461) => x"00", (0 + 6462) => x"00", (0 + 6463) => x"00", (0 + 6464) => x"00", (0 + 6465) => x"00", (0 + 6466) => x"00", (0 + 6467) => x"00", (0 + 6468) => x"00", (0 + 6469) => x"00", (0 + 6470) => x"00", (0 + 6471) => x"00", (0 + 6472) => x"00", (0 + 6473) => x"00", (0 + 6474) => x"00", (0 + 6475) => x"00", (0 + 6476) => x"00", (0 + 6477) => x"00", (0 + 6478) => x"00", (0 + 6479) => x"00", (0 + 6480) => x"00", (0 + 6481) => x"00", (0 + 6482) => x"00", (0 + 6483) => x"00", (0 + 6484) => x"00", (0 + 6485) => x"00", (0 + 6486) => x"00", (0 + 6487) => x"00", (0 + 6488) => x"00", (0 + 6489) => x"00", (0 + 6490) => x"00", (0 + 6491) => x"00", (0 + 6492) => x"00", (0 + 6493) => x"00", (0 + 6494) => x"00", (0 + 6495) => x"00", (0 + 6496) => x"00", (0 + 6497) => x"00", (0 + 6498) => x"00", (0 + 6499) => x"00", (0 + 6500) => x"00", (0 + 6501) => x"00", (0 + 6502) => x"00", (0 + 6503) => x"00", (0 + 6504) => x"00", (0 + 6505) => x"00", (0 + 6506) => x"00", (0 + 6507) => x"00", (0 + 6508) => x"00", (0 + 6509) => x"00", (0 + 6510) => x"00", (0 + 6511) => x"00", (0 + 6512) => x"00", (0 + 6513) => x"00", (0 + 6514) => x"00", (0 + 6515) => x"00", (0 + 6516) => x"00", (0 + 6517) => x"00", (0 + 6518) => x"00", (0 + 6519) => x"00", (0 + 6520) => x"00", (0 + 6521) => x"00", (0 + 6522) => x"00", (0 + 6523) => x"00", (0 + 6524) => x"00", (0 + 6525) => x"00", (0 + 6526) => x"00", (0 + 6527) => x"00", (0 + 6528) => x"00", (0 + 6529) => x"00", (0 + 6530) => x"00", (0 + 6531) => x"00", (0 + 6532) => x"00", (0 + 6533) => x"00", (0 + 6534) => x"00", (0 + 6535) => x"00", (0 + 6536) => x"00", (0 + 6537) => x"00", (0 + 6538) => x"00", (0 + 6539) => x"00", (0 + 6540) => x"00", (0 + 6541) => x"00", (0 + 6542) => x"00", (0 + 6543) => x"00", (0 + 6544) => x"00", (0 + 6545) => x"00", (0 + 6546) => x"00", (0 + 6547) => x"00", (0 + 6548) => x"00", (0 + 6549) => x"00", (0 + 6550) => x"00", (0 + 6551) => x"00", (0 + 6552) => x"00", (0 + 6553) => x"00", (0 + 6554) => x"00", (0 + 6555) => x"00", (0 + 6556) => x"00", (0 + 6557) => x"00", (0 + 6558) => x"00", (0 + 6559) => x"00", (0 + 6560) => x"00", (0 + 6561) => x"00", (0 + 6562) => x"00", (0 + 6563) => x"00", (0 + 6564) => x"00", (0 + 6565) => x"00", (0 + 6566) => x"00", (0 + 6567) => x"00", (0 + 6568) => x"00", (0 + 6569) => x"00", (0 + 6570) => x"00", (0 + 6571) => x"00", (0 + 6572) => x"00", (0 + 6573) => x"00", (0 + 6574) => x"00", (0 + 6575) => x"00", (0 + 6576) => x"00", (0 + 6577) => x"00", (0 + 6578) => x"00", (0 + 6579) => x"00", (0 + 6580) => x"00", (0 + 6581) => x"00", (0 + 6582) => x"00", (0 + 6583) => x"00", (0 + 6584) => x"00", (0 + 6585) => x"00", (0 + 6586) => x"00", (0 + 6587) => x"00", (0 + 6588) => x"00", (0 + 6589) => x"00", (0 + 6590) => x"00", (0 + 6591) => x"00", (0 + 6592) => x"00", (0 + 6593) => x"00", (0 + 6594) => x"00", (0 + 6595) => x"00", (0 + 6596) => x"00", (0 + 6597) => x"00", (0 + 6598) => x"00", (0 + 6599) => x"00", (0 + 6600) => x"00", (0 + 6601) => x"00", (0 + 6602) => x"00", (0 + 6603) => x"00", (0 + 6604) => x"00", (0 + 6605) => x"00", (0 + 6606) => x"00", (0 + 6607) => x"00", (0 + 6608) => x"00", (0 + 6609) => x"00", (0 + 6610) => x"00", (0 + 6611) => x"00", (0 + 6612) => x"00", (0 + 6613) => x"00", (0 + 6614) => x"00", (0 + 6615) => x"00", (0 + 6616) => x"00", (0 + 6617) => x"00", (0 + 6618) => x"00", (0 + 6619) => x"00", (0 + 6620) => x"00", (0 + 6621) => x"00", (0 + 6622) => x"00", (0 + 6623) => x"00", (0 + 6624) => x"00", (0 + 6625) => x"00", (0 + 6626) => x"00", (0 + 6627) => x"00", (0 + 6628) => x"00", (0 + 6629) => x"00", (0 + 6630) => x"00", (0 + 6631) => x"00", (0 + 6632) => x"00", (0 + 6633) => x"00", (0 + 6634) => x"00", (0 + 6635) => x"00", (0 + 6636) => x"00", (0 + 6637) => x"00", (0 + 6638) => x"00", (0 + 6639) => x"00", (0 + 6640) => x"00", (0 + 6641) => x"00", (0 + 6642) => x"00", (0 + 6643) => x"00", (0 + 6644) => x"00", (0 + 6645) => x"00", (0 + 6646) => x"00", (0 + 6647) => x"00", (0 + 6648) => x"00", (0 + 6649) => x"00", (0 + 6650) => x"00", (0 + 6651) => x"00", (0 + 6652) => x"00", (0 + 6653) => x"00", (0 + 6654) => x"00", (0 + 6655) => x"00", (0 + 6656) => x"00", (0 + 6657) => x"00", (0 + 6658) => x"00", (0 + 6659) => x"00", (0 + 6660) => x"00", (0 + 6661) => x"00", (0 + 6662) => x"00", (0 + 6663) => x"00", (0 + 6664) => x"00", (0 + 6665) => x"00", (0 + 6666) => x"00", (0 + 6667) => x"00", (0 + 6668) => x"00", (0 + 6669) => x"00", (0 + 6670) => x"00", (0 + 6671) => x"00", (0 + 6672) => x"00", (0 + 6673) => x"00", (0 + 6674) => x"00", (0 + 6675) => x"00", (0 + 6676) => x"00", (0 + 6677) => x"00", (0 + 6678) => x"00", (0 + 6679) => x"00", (0 + 6680) => x"00", (0 + 6681) => x"00", (0 + 6682) => x"00", (0 + 6683) => x"00", (0 + 6684) => x"00", (0 + 6685) => x"00", (0 + 6686) => x"00", (0 + 6687) => x"00", (0 + 6688) => x"00", (0 + 6689) => x"00", (0 + 6690) => x"00", (0 + 6691) => x"00", (0 + 6692) => x"00", (0 + 6693) => x"00", (0 + 6694) => x"00", (0 + 6695) => x"00", (0 + 6696) => x"00", (0 + 6697) => x"00", (0 + 6698) => x"00", (0 + 6699) => x"00", (0 + 6700) => x"00", (0 + 6701) => x"00", (0 + 6702) => x"00", (0 + 6703) => x"00", (0 + 6704) => x"00", (0 + 6705) => x"00", (0 + 6706) => x"00", (0 + 6707) => x"00", (0 + 6708) => x"00", (0 + 6709) => x"00", (0 + 6710) => x"00", (0 + 6711) => x"00", (0 + 6712) => x"00", (0 + 6713) => x"00", (0 + 6714) => x"00", (0 + 6715) => x"00", (0 + 6716) => x"00", (0 + 6717) => x"00", (0 + 6718) => x"00", (0 + 6719) => x"00", (0 + 6720) => x"00", (0 + 6721) => x"00", (0 + 6722) => x"00", (0 + 6723) => x"00", (0 + 6724) => x"00", (0 + 6725) => x"00", (0 + 6726) => x"00", (0 + 6727) => x"00", (0 + 6728) => x"00", (0 + 6729) => x"00", (0 + 6730) => x"00", (0 + 6731) => x"00", (0 + 6732) => x"00", (0 + 6733) => x"00", (0 + 6734) => x"00", (0 + 6735) => x"00", (0 + 6736) => x"00", (0 + 6737) => x"00", (0 + 6738) => x"00", (0 + 6739) => x"00", (0 + 6740) => x"00", (0 + 6741) => x"00", (0 + 6742) => x"00", (0 + 6743) => x"00", (0 + 6744) => x"00", (0 + 6745) => x"00", (0 + 6746) => x"00", (0 + 6747) => x"00", (0 + 6748) => x"00", (0 + 6749) => x"00", (0 + 6750) => x"00", (0 + 6751) => x"00", (0 + 6752) => x"00", (0 + 6753) => x"00", (0 + 6754) => x"00", (0 + 6755) => x"00", (0 + 6756) => x"00", (0 + 6757) => x"00", (0 + 6758) => x"00", (0 + 6759) => x"00", (0 + 6760) => x"00", (0 + 6761) => x"00", (0 + 6762) => x"00", (0 + 6763) => x"00", (0 + 6764) => x"00", (0 + 6765) => x"00", (0 + 6766) => x"00", (0 + 6767) => x"00", (0 + 6768) => x"00", (0 + 6769) => x"00", (0 + 6770) => x"00", (0 + 6771) => x"00", (0 + 6772) => x"00", (0 + 6773) => x"00", (0 + 6774) => x"00", (0 + 6775) => x"00", (0 + 6776) => x"00", (0 + 6777) => x"00", (0 + 6778) => x"00", (0 + 6779) => x"00", (0 + 6780) => x"00", (0 + 6781) => x"00", (0 + 6782) => x"00", (0 + 6783) => x"00", (0 + 6784) => x"00", (0 + 6785) => x"00", (0 + 6786) => x"00", (0 + 6787) => x"00", (0 + 6788) => x"00", (0 + 6789) => x"00", (0 + 6790) => x"00", (0 + 6791) => x"00", (0 + 6792) => x"00", (0 + 6793) => x"00", (0 + 6794) => x"00", (0 + 6795) => x"00", (0 + 6796) => x"00", (0 + 6797) => x"00", (0 + 6798) => x"00", (0 + 6799) => x"00", (0 + 6800) => x"00", (0 + 6801) => x"00", (0 + 6802) => x"00", (0 + 6803) => x"00", (0 + 6804) => x"00", (0 + 6805) => x"00", (0 + 6806) => x"00", (0 + 6807) => x"00", (0 + 6808) => x"00", (0 + 6809) => x"00", (0 + 6810) => x"00", (0 + 6811) => x"00", (0 + 6812) => x"00", (0 + 6813) => x"00", (0 + 6814) => x"00", (0 + 6815) => x"00", (0 + 6816) => x"00", (0 + 6817) => x"00", (0 + 6818) => x"00", (0 + 6819) => x"00", (0 + 6820) => x"00", (0 + 6821) => x"00", (0 + 6822) => x"00", (0 + 6823) => x"00", (0 + 6824) => x"00", (0 + 6825) => x"00", (0 + 6826) => x"00", (0 + 6827) => x"00", (0 + 6828) => x"00", (0 + 6829) => x"00", (0 + 6830) => x"00", (0 + 6831) => x"00", (0 + 6832) => x"00", (0 + 6833) => x"00", (0 + 6834) => x"00", (0 + 6835) => x"00", (0 + 6836) => x"00", (0 + 6837) => x"00", (0 + 6838) => x"00", (0 + 6839) => x"00", (0 + 6840) => x"00", (0 + 6841) => x"00", (0 + 6842) => x"00", (0 + 6843) => x"00", (0 + 6844) => x"00", (0 + 6845) => x"00", (0 + 6846) => x"00", (0 + 6847) => x"00", (0 + 6848) => x"00", (0 + 6849) => x"00", (0 + 6850) => x"00", (0 + 6851) => x"00", (0 + 6852) => x"00", (0 + 6853) => x"00", (0 + 6854) => x"00", (0 + 6855) => x"00", (0 + 6856) => x"00", (0 + 6857) => x"00", (0 + 6858) => x"00", (0 + 6859) => x"00", (0 + 6860) => x"00", (0 + 6861) => x"00", (0 + 6862) => x"00", (0 + 6863) => x"00", (0 + 6864) => x"00", (0 + 6865) => x"00", (0 + 6866) => x"00", (0 + 6867) => x"00", (0 + 6868) => x"00", (0 + 6869) => x"00", (0 + 6870) => x"00", (0 + 6871) => x"00", (0 + 6872) => x"00", (0 + 6873) => x"00", (0 + 6874) => x"00", (0 + 6875) => x"00", (0 + 6876) => x"00", (0 + 6877) => x"00", (0 + 6878) => x"00", (0 + 6879) => x"00", (0 + 6880) => x"00", (0 + 6881) => x"00", (0 + 6882) => x"00", (0 + 6883) => x"00", (0 + 6884) => x"00", (0 + 6885) => x"00", (0 + 6886) => x"00", (0 + 6887) => x"00", (0 + 6888) => x"00", (0 + 6889) => x"00", (0 + 6890) => x"00", (0 + 6891) => x"00", (0 + 6892) => x"00", (0 + 6893) => x"00", (0 + 6894) => x"00", (0 + 6895) => x"00", (0 + 6896) => x"00", (0 + 6897) => x"00", (0 + 6898) => x"00", (0 + 6899) => x"00", (0 + 6900) => x"00", (0 + 6901) => x"00", (0 + 6902) => x"00", (0 + 6903) => x"00", (0 + 6904) => x"00", (0 + 6905) => x"00", (0 + 6906) => x"00", (0 + 6907) => x"00", (0 + 6908) => x"00", (0 + 6909) => x"00", (0 + 6910) => x"00", (0 + 6911) => x"00", (0 + 6912) => x"00", (0 + 6913) => x"00", (0 + 6914) => x"00", (0 + 6915) => x"00", (0 + 6916) => x"00", (0 + 6917) => x"00", (0 + 6918) => x"00", (0 + 6919) => x"00", (0 + 6920) => x"00", (0 + 6921) => x"00", (0 + 6922) => x"00", (0 + 6923) => x"00", (0 + 6924) => x"00", (0 + 6925) => x"00", (0 + 6926) => x"00", (0 + 6927) => x"00", (0 + 6928) => x"00", (0 + 6929) => x"00", (0 + 6930) => x"00", (0 + 6931) => x"00", (0 + 6932) => x"00", (0 + 6933) => x"00", (0 + 6934) => x"00", (0 + 6935) => x"00", (0 + 6936) => x"00", (0 + 6937) => x"00", (0 + 6938) => x"00", (0 + 6939) => x"00", (0 + 6940) => x"00", (0 + 6941) => x"00", (0 + 6942) => x"00", (0 + 6943) => x"00", (0 + 6944) => x"00", (0 + 6945) => x"00", (0 + 6946) => x"00", (0 + 6947) => x"00", (0 + 6948) => x"00", (0 + 6949) => x"00", (0 + 6950) => x"00", (0 + 6951) => x"00", (0 + 6952) => x"00", (0 + 6953) => x"00", (0 + 6954) => x"00", (0 + 6955) => x"00", (0 + 6956) => x"00", (0 + 6957) => x"00", (0 + 6958) => x"00", (0 + 6959) => x"00", (0 + 6960) => x"00", (0 + 6961) => x"00", (0 + 6962) => x"00", (0 + 6963) => x"00", (0 + 6964) => x"00", (0 + 6965) => x"00", (0 + 6966) => x"00", (0 + 6967) => x"00", (0 + 6968) => x"00", (0 + 6969) => x"00", (0 + 6970) => x"00", (0 + 6971) => x"00", (0 + 6972) => x"00", (0 + 6973) => x"00", (0 + 6974) => x"00", (0 + 6975) => x"00", (0 + 6976) => x"00", (0 + 6977) => x"00", (0 + 6978) => x"00", (0 + 6979) => x"00", (0 + 6980) => x"00", (0 + 6981) => x"00", (0 + 6982) => x"00", (0 + 6983) => x"00", (0 + 6984) => x"00", (0 + 6985) => x"00", (0 + 6986) => x"00", (0 + 6987) => x"00", (0 + 6988) => x"00", (0 + 6989) => x"00", (0 + 6990) => x"00", (0 + 6991) => x"00", (0 + 6992) => x"00", (0 + 6993) => x"00", (0 + 6994) => x"00", (0 + 6995) => x"00", (0 + 6996) => x"00", (0 + 6997) => x"00", (0 + 6998) => x"00", (0 + 6999) => x"00", (0 + 7000) => x"00", (0 + 7001) => x"00", (0 + 7002) => x"00", (0 + 7003) => x"00", (0 + 7004) => x"00", (0 + 7005) => x"00", (0 + 7006) => x"00", (0 + 7007) => x"00", (0 + 7008) => x"00", (0 + 7009) => x"00", (0 + 7010) => x"00", (0 + 7011) => x"00", (0 + 7012) => x"00", (0 + 7013) => x"00", (0 + 7014) => x"00", (0 + 7015) => x"00", (0 + 7016) => x"00", (0 + 7017) => x"00", (0 + 7018) => x"00", (0 + 7019) => x"00", (0 + 7020) => x"00", (0 + 7021) => x"00", (0 + 7022) => x"00", (0 + 7023) => x"00", (0 + 7024) => x"00", (0 + 7025) => x"00", (0 + 7026) => x"00", (0 + 7027) => x"00", (0 + 7028) => x"00", (0 + 7029) => x"00", (0 + 7030) => x"00", (0 + 7031) => x"00", (0 + 7032) => x"00", (0 + 7033) => x"00", (0 + 7034) => x"00", (0 + 7035) => x"00", (0 + 7036) => x"00", (0 + 7037) => x"00", (0 + 7038) => x"00", (0 + 7039) => x"00", (0 + 7040) => x"00", (0 + 7041) => x"00", (0 + 7042) => x"00", (0 + 7043) => x"00", (0 + 7044) => x"00", (0 + 7045) => x"00", (0 + 7046) => x"00", (0 + 7047) => x"00", (0 + 7048) => x"00", (0 + 7049) => x"00", (0 + 7050) => x"00", (0 + 7051) => x"00", (0 + 7052) => x"00", (0 + 7053) => x"00", (0 + 7054) => x"00", (0 + 7055) => x"00", (0 + 7056) => x"00", (0 + 7057) => x"00", (0 + 7058) => x"00", (0 + 7059) => x"00", (0 + 7060) => x"00", (0 + 7061) => x"00", (0 + 7062) => x"00", (0 + 7063) => x"00", (0 + 7064) => x"00", (0 + 7065) => x"00", (0 + 7066) => x"00", (0 + 7067) => x"00", (0 + 7068) => x"00", (0 + 7069) => x"00", (0 + 7070) => x"00", (0 + 7071) => x"00", (0 + 7072) => x"00", (0 + 7073) => x"00", (0 + 7074) => x"00", (0 + 7075) => x"00", (0 + 7076) => x"00", (0 + 7077) => x"00", (0 + 7078) => x"00", (0 + 7079) => x"00", (0 + 7080) => x"00", (0 + 7081) => x"00", (0 + 7082) => x"00", (0 + 7083) => x"00", (0 + 7084) => x"00", (0 + 7085) => x"00", (0 + 7086) => x"00", (0 + 7087) => x"00", (0 + 7088) => x"00", (0 + 7089) => x"00", (0 + 7090) => x"00", (0 + 7091) => x"00", (0 + 7092) => x"00", (0 + 7093) => x"00", (0 + 7094) => x"00", (0 + 7095) => x"00", (0 + 7096) => x"00", (0 + 7097) => x"00", (0 + 7098) => x"00", (0 + 7099) => x"00", (0 + 7100) => x"00", (0 + 7101) => x"00", (0 + 7102) => x"00", (0 + 7103) => x"00", (0 + 7104) => x"00", (0 + 7105) => x"00", (0 + 7106) => x"00", (0 + 7107) => x"00", (0 + 7108) => x"00", (0 + 7109) => x"00", (0 + 7110) => x"00", (0 + 7111) => x"00", (0 + 7112) => x"00", (0 + 7113) => x"00", (0 + 7114) => x"00", (0 + 7115) => x"00", (0 + 7116) => x"00", (0 + 7117) => x"00", (0 + 7118) => x"00", (0 + 7119) => x"00", (0 + 7120) => x"00", (0 + 7121) => x"00", (0 + 7122) => x"00", (0 + 7123) => x"00", (0 + 7124) => x"00", (0 + 7125) => x"00", (0 + 7126) => x"00", (0 + 7127) => x"00", (0 + 7128) => x"00", (0 + 7129) => x"00", (0 + 7130) => x"00", (0 + 7131) => x"00", (0 + 7132) => x"00", (0 + 7133) => x"00", (0 + 7134) => x"00", (0 + 7135) => x"00", (0 + 7136) => x"00", (0 + 7137) => x"00", (0 + 7138) => x"00", (0 + 7139) => x"00", (0 + 7140) => x"00", (0 + 7141) => x"00", (0 + 7142) => x"00", (0 + 7143) => x"00", (0 + 7144) => x"00", (0 + 7145) => x"00", (0 + 7146) => x"00", (0 + 7147) => x"00", (0 + 7148) => x"00", (0 + 7149) => x"00", (0 + 7150) => x"00", (0 + 7151) => x"00", (0 + 7152) => x"00", (0 + 7153) => x"00", (0 + 7154) => x"00", (0 + 7155) => x"00", (0 + 7156) => x"00", (0 + 7157) => x"00", (0 + 7158) => x"00", (0 + 7159) => x"00", (0 + 7160) => x"00", (0 + 7161) => x"00", (0 + 7162) => x"00", (0 + 7163) => x"00", (0 + 7164) => x"00", (0 + 7165) => x"00", (0 + 7166) => x"00", (0 + 7167) => x"00", (0 + 7168) => x"00", (0 + 7169) => x"00", (0 + 7170) => x"00", (0 + 7171) => x"00", (0 + 7172) => x"00", (0 + 7173) => x"00", (0 + 7174) => x"00", (0 + 7175) => x"00", (0 + 7176) => x"00", (0 + 7177) => x"00", (0 + 7178) => x"00", (0 + 7179) => x"00", (0 + 7180) => x"00", (0 + 7181) => x"00", (0 + 7182) => x"00", (0 + 7183) => x"00", (0 + 7184) => x"00", (0 + 7185) => x"00", (0 + 7186) => x"00", (0 + 7187) => x"00", (0 + 7188) => x"00", (0 + 7189) => x"00", (0 + 7190) => x"00", (0 + 7191) => x"00", (0 + 7192) => x"00", (0 + 7193) => x"00", (0 + 7194) => x"00", (0 + 7195) => x"00", (0 + 7196) => x"00", (0 + 7197) => x"00", (0 + 7198) => x"00", (0 + 7199) => x"00", (0 + 7200) => x"00", (0 + 7201) => x"00", (0 + 7202) => x"00", (0 + 7203) => x"00", (0 + 7204) => x"00", (0 + 7205) => x"00", (0 + 7206) => x"00", (0 + 7207) => x"00", (0 + 7208) => x"00", (0 + 7209) => x"00", (0 + 7210) => x"00", (0 + 7211) => x"00", (0 + 7212) => x"00", (0 + 7213) => x"00", (0 + 7214) => x"00", (0 + 7215) => x"00", (0 + 7216) => x"00", (0 + 7217) => x"00", (0 + 7218) => x"00", (0 + 7219) => x"00", (0 + 7220) => x"00", (0 + 7221) => x"00", (0 + 7222) => x"00", (0 + 7223) => x"00", (0 + 7224) => x"00", (0 + 7225) => x"00", (0 + 7226) => x"00", (0 + 7227) => x"00", (0 + 7228) => x"00", (0 + 7229) => x"00", (0 + 7230) => x"00", (0 + 7231) => x"00", (0 + 7232) => x"00", (0 + 7233) => x"00", (0 + 7234) => x"00", (0 + 7235) => x"00", (0 + 7236) => x"00", (0 + 7237) => x"00", (0 + 7238) => x"00", (0 + 7239) => x"00", (0 + 7240) => x"00", (0 + 7241) => x"00", (0 + 7242) => x"00", (0 + 7243) => x"00", (0 + 7244) => x"00", (0 + 7245) => x"00", (0 + 7246) => x"00", (0 + 7247) => x"00", (0 + 7248) => x"00", (0 + 7249) => x"00", (0 + 7250) => x"00", (0 + 7251) => x"00", (0 + 7252) => x"00", (0 + 7253) => x"00", (0 + 7254) => x"00", (0 + 7255) => x"00", (0 + 7256) => x"00", (0 + 7257) => x"00", (0 + 7258) => x"00", (0 + 7259) => x"00", (0 + 7260) => x"00", (0 + 7261) => x"00", (0 + 7262) => x"00", (0 + 7263) => x"00", (0 + 7264) => x"00", (0 + 7265) => x"00", (0 + 7266) => x"00", (0 + 7267) => x"00", (0 + 7268) => x"00", (0 + 7269) => x"00", (0 + 7270) => x"00", (0 + 7271) => x"00", (0 + 7272) => x"00", (0 + 7273) => x"00", (0 + 7274) => x"00", (0 + 7275) => x"00", (0 + 7276) => x"00", (0 + 7277) => x"00", (0 + 7278) => x"00", (0 + 7279) => x"00", (0 + 7280) => x"00", (0 + 7281) => x"00", (0 + 7282) => x"00", (0 + 7283) => x"00", (0 + 7284) => x"00", (0 + 7285) => x"00", (0 + 7286) => x"00", (0 + 7287) => x"00", (0 + 7288) => x"00", (0 + 7289) => x"00", (0 + 7290) => x"00", (0 + 7291) => x"00", (0 + 7292) => x"00", (0 + 7293) => x"00", (0 + 7294) => x"00", (0 + 7295) => x"00", (0 + 7296) => x"00", (0 + 7297) => x"00", (0 + 7298) => x"00", (0 + 7299) => x"00", (0 + 7300) => x"00", (0 + 7301) => x"00", (0 + 7302) => x"00", (0 + 7303) => x"00", (0 + 7304) => x"00", (0 + 7305) => x"00", (0 + 7306) => x"00", (0 + 7307) => x"00", (0 + 7308) => x"00", (0 + 7309) => x"00", (0 + 7310) => x"00", (0 + 7311) => x"00", (0 + 7312) => x"00", (0 + 7313) => x"00", (0 + 7314) => x"00", (0 + 7315) => x"00", (0 + 7316) => x"00", (0 + 7317) => x"00", (0 + 7318) => x"00", (0 + 7319) => x"00", (0 + 7320) => x"00", (0 + 7321) => x"00", (0 + 7322) => x"00", (0 + 7323) => x"00", (0 + 7324) => x"00", (0 + 7325) => x"00", (0 + 7326) => x"00", (0 + 7327) => x"00", (0 + 7328) => x"00", (0 + 7329) => x"00", (0 + 7330) => x"00", (0 + 7331) => x"00", (0 + 7332) => x"00", (0 + 7333) => x"00", (0 + 7334) => x"00", (0 + 7335) => x"00", (0 + 7336) => x"00", (0 + 7337) => x"00", (0 + 7338) => x"00", (0 + 7339) => x"00", (0 + 7340) => x"00", (0 + 7341) => x"00", (0 + 7342) => x"00", (0 + 7343) => x"00", (0 + 7344) => x"00", (0 + 7345) => x"00", (0 + 7346) => x"00", (0 + 7347) => x"00", (0 + 7348) => x"00", (0 + 7349) => x"00", (0 + 7350) => x"00", (0 + 7351) => x"00", (0 + 7352) => x"00", (0 + 7353) => x"00", (0 + 7354) => x"00", (0 + 7355) => x"00", (0 + 7356) => x"00", (0 + 7357) => x"00", (0 + 7358) => x"00", (0 + 7359) => x"00", (0 + 7360) => x"00", (0 + 7361) => x"00", (0 + 7362) => x"00", (0 + 7363) => x"00", (0 + 7364) => x"00", (0 + 7365) => x"00", (0 + 7366) => x"00", (0 + 7367) => x"00", (0 + 7368) => x"00", (0 + 7369) => x"00", (0 + 7370) => x"00", (0 + 7371) => x"00", (0 + 7372) => x"00", (0 + 7373) => x"00", (0 + 7374) => x"00", (0 + 7375) => x"00", (0 + 7376) => x"00", (0 + 7377) => x"00", (0 + 7378) => x"00", (0 + 7379) => x"00", (0 + 7380) => x"00", (0 + 7381) => x"00", (0 + 7382) => x"00", (0 + 7383) => x"00", (0 + 7384) => x"00", (0 + 7385) => x"00", (0 + 7386) => x"00", (0 + 7387) => x"00", (0 + 7388) => x"00", (0 + 7389) => x"00", (0 + 7390) => x"00", (0 + 7391) => x"00", (0 + 7392) => x"00", (0 + 7393) => x"00", (0 + 7394) => x"00", (0 + 7395) => x"00", (0 + 7396) => x"00", (0 + 7397) => x"00", (0 + 7398) => x"00", (0 + 7399) => x"00", (0 + 7400) => x"00", (0 + 7401) => x"00", (0 + 7402) => x"00", (0 + 7403) => x"00", (0 + 7404) => x"00", (0 + 7405) => x"00", (0 + 7406) => x"00", (0 + 7407) => x"00", (0 + 7408) => x"00", (0 + 7409) => x"00", (0 + 7410) => x"00", (0 + 7411) => x"00", (0 + 7412) => x"00", (0 + 7413) => x"00", (0 + 7414) => x"00", (0 + 7415) => x"00", (0 + 7416) => x"00", (0 + 7417) => x"00", (0 + 7418) => x"00", (0 + 7419) => x"00", (0 + 7420) => x"00", (0 + 7421) => x"00", (0 + 7422) => x"00", (0 + 7423) => x"00", (0 + 7424) => x"00", (0 + 7425) => x"00", (0 + 7426) => x"00", (0 + 7427) => x"00", (0 + 7428) => x"00", (0 + 7429) => x"00", (0 + 7430) => x"00", (0 + 7431) => x"00", (0 + 7432) => x"00", (0 + 7433) => x"00", (0 + 7434) => x"00", (0 + 7435) => x"00", (0 + 7436) => x"00", (0 + 7437) => x"00", (0 + 7438) => x"00", (0 + 7439) => x"00", (0 + 7440) => x"00", (0 + 7441) => x"00", (0 + 7442) => x"00", (0 + 7443) => x"00", (0 + 7444) => x"00", (0 + 7445) => x"00", (0 + 7446) => x"00", (0 + 7447) => x"00", (0 + 7448) => x"00", (0 + 7449) => x"00", (0 + 7450) => x"00", (0 + 7451) => x"00", (0 + 7452) => x"00", (0 + 7453) => x"00", (0 + 7454) => x"00", (0 + 7455) => x"00", (0 + 7456) => x"00", (0 + 7457) => x"00", (0 + 7458) => x"00", (0 + 7459) => x"00", (0 + 7460) => x"00", (0 + 7461) => x"00", (0 + 7462) => x"00", (0 + 7463) => x"00", (0 + 7464) => x"00", (0 + 7465) => x"00", (0 + 7466) => x"00", (0 + 7467) => x"00", (0 + 7468) => x"00", (0 + 7469) => x"00", (0 + 7470) => x"00", (0 + 7471) => x"00", (0 + 7472) => x"00", (0 + 7473) => x"00", (0 + 7474) => x"00", (0 + 7475) => x"00", (0 + 7476) => x"00", (0 + 7477) => x"00", (0 + 7478) => x"00", (0 + 7479) => x"00", (0 + 7480) => x"00", (0 + 7481) => x"00", (0 + 7482) => x"00", (0 + 7483) => x"00", (0 + 7484) => x"00", (0 + 7485) => x"00", (0 + 7486) => x"00", (0 + 7487) => x"00", (0 + 7488) => x"00", (0 + 7489) => x"00", (0 + 7490) => x"00", (0 + 7491) => x"00", (0 + 7492) => x"00", (0 + 7493) => x"00", (0 + 7494) => x"00", (0 + 7495) => x"00", (0 + 7496) => x"00", (0 + 7497) => x"00", (0 + 7498) => x"00", (0 + 7499) => x"00", (0 + 7500) => x"00", (0 + 7501) => x"00", (0 + 7502) => x"00", (0 + 7503) => x"00", (0 + 7504) => x"00", (0 + 7505) => x"00", (0 + 7506) => x"00", (0 + 7507) => x"00", (0 + 7508) => x"00", (0 + 7509) => x"00", (0 + 7510) => x"00", (0 + 7511) => x"00", (0 + 7512) => x"00", (0 + 7513) => x"00", (0 + 7514) => x"00", (0 + 7515) => x"00", (0 + 7516) => x"00", (0 + 7517) => x"00", (0 + 7518) => x"00", (0 + 7519) => x"00", (0 + 7520) => x"00", (0 + 7521) => x"00", (0 + 7522) => x"00", (0 + 7523) => x"00", (0 + 7524) => x"00", (0 + 7525) => x"00", (0 + 7526) => x"00", (0 + 7527) => x"00", (0 + 7528) => x"00", (0 + 7529) => x"00", (0 + 7530) => x"00", (0 + 7531) => x"00", (0 + 7532) => x"00", (0 + 7533) => x"00", (0 + 7534) => x"00", (0 + 7535) => x"00", (0 + 7536) => x"00", (0 + 7537) => x"00", (0 + 7538) => x"00", (0 + 7539) => x"00", (0 + 7540) => x"00", (0 + 7541) => x"00", (0 + 7542) => x"00", (0 + 7543) => x"00", (0 + 7544) => x"00", (0 + 7545) => x"00", (0 + 7546) => x"00", (0 + 7547) => x"00", (0 + 7548) => x"00", (0 + 7549) => x"00", (0 + 7550) => x"00", (0 + 7551) => x"00", (0 + 7552) => x"00", (0 + 7553) => x"00", (0 + 7554) => x"00", (0 + 7555) => x"00", (0 + 7556) => x"00", (0 + 7557) => x"00", (0 + 7558) => x"00", (0 + 7559) => x"00", (0 + 7560) => x"00", (0 + 7561) => x"00", (0 + 7562) => x"00", (0 + 7563) => x"00", (0 + 7564) => x"00", (0 + 7565) => x"00", (0 + 7566) => x"00", (0 + 7567) => x"00", (0 + 7568) => x"00", (0 + 7569) => x"00", (0 + 7570) => x"00", (0 + 7571) => x"00", (0 + 7572) => x"00", (0 + 7573) => x"00", (0 + 7574) => x"00", (0 + 7575) => x"00", (0 + 7576) => x"00", (0 + 7577) => x"00", (0 + 7578) => x"00", (0 + 7579) => x"00", (0 + 7580) => x"00", (0 + 7581) => x"00", (0 + 7582) => x"00", (0 + 7583) => x"00", (0 + 7584) => x"00", (0 + 7585) => x"00", (0 + 7586) => x"00", (0 + 7587) => x"00", (0 + 7588) => x"00", (0 + 7589) => x"00", (0 + 7590) => x"00", (0 + 7591) => x"00", (0 + 7592) => x"00", (0 + 7593) => x"00", (0 + 7594) => x"00", (0 + 7595) => x"00", (0 + 7596) => x"00", (0 + 7597) => x"00", (0 + 7598) => x"00", (0 + 7599) => x"00", (0 + 7600) => x"00", (0 + 7601) => x"00", (0 + 7602) => x"00", (0 + 7603) => x"00", (0 + 7604) => x"00", (0 + 7605) => x"00", (0 + 7606) => x"00", (0 + 7607) => x"00", (0 + 7608) => x"00", (0 + 7609) => x"00", (0 + 7610) => x"00", (0 + 7611) => x"00", (0 + 7612) => x"00", (0 + 7613) => x"00", (0 + 7614) => x"00", (0 + 7615) => x"00", (0 + 7616) => x"00", (0 + 7617) => x"00", (0 + 7618) => x"00", (0 + 7619) => x"00", (0 + 7620) => x"00", (0 + 7621) => x"00", (0 + 7622) => x"00", (0 + 7623) => x"00", (0 + 7624) => x"00", (0 + 7625) => x"00", (0 + 7626) => x"00", (0 + 7627) => x"00", (0 + 7628) => x"00", (0 + 7629) => x"00", (0 + 7630) => x"00", (0 + 7631) => x"00", (0 + 7632) => x"00", (0 + 7633) => x"00", (0 + 7634) => x"00", (0 + 7635) => x"00", (0 + 7636) => x"00", (0 + 7637) => x"00", (0 + 7638) => x"00", (0 + 7639) => x"00", (0 + 7640) => x"00", (0 + 7641) => x"00", (0 + 7642) => x"00", (0 + 7643) => x"00", (0 + 7644) => x"00", (0 + 7645) => x"00", (0 + 7646) => x"00", (0 + 7647) => x"00", (0 + 7648) => x"00", (0 + 7649) => x"00", (0 + 7650) => x"00", (0 + 7651) => x"00", (0 + 7652) => x"00", (0 + 7653) => x"00", (0 + 7654) => x"00", (0 + 7655) => x"00", (0 + 7656) => x"00", (0 + 7657) => x"00", (0 + 7658) => x"00", (0 + 7659) => x"00", (0 + 7660) => x"00", (0 + 7661) => x"00", (0 + 7662) => x"00", (0 + 7663) => x"00", (0 + 7664) => x"00", (0 + 7665) => x"00", (0 + 7666) => x"00", (0 + 7667) => x"00", (0 + 7668) => x"00", (0 + 7669) => x"00", (0 + 7670) => x"00", (0 + 7671) => x"00", (0 + 7672) => x"00", (0 + 7673) => x"00", (0 + 7674) => x"00", (0 + 7675) => x"00", (0 + 7676) => x"00", (0 + 7677) => x"00", (0 + 7678) => x"00", (0 + 7679) => x"00", (0 + 7680) => x"00", (0 + 7681) => x"00", (0 + 7682) => x"00", (0 + 7683) => x"00", (0 + 7684) => x"00", (0 + 7685) => x"00", (0 + 7686) => x"00", (0 + 7687) => x"00", (0 + 7688) => x"00", (0 + 7689) => x"00", (0 + 7690) => x"00", (0 + 7691) => x"00", (0 + 7692) => x"00", (0 + 7693) => x"00", (0 + 7694) => x"00", (0 + 7695) => x"00", (0 + 7696) => x"00", (0 + 7697) => x"00", (0 + 7698) => x"00", (0 + 7699) => x"00", (0 + 7700) => x"00", (0 + 7701) => x"00", (0 + 7702) => x"00", (0 + 7703) => x"00", (0 + 7704) => x"00", (0 + 7705) => x"00", (0 + 7706) => x"00", (0 + 7707) => x"00", (0 + 7708) => x"00", (0 + 7709) => x"00", (0 + 7710) => x"00", (0 + 7711) => x"00", (0 + 7712) => x"00", (0 + 7713) => x"00", (0 + 7714) => x"00", (0 + 7715) => x"00", (0 + 7716) => x"00", (0 + 7717) => x"00", (0 + 7718) => x"00", (0 + 7719) => x"00", (0 + 7720) => x"00", (0 + 7721) => x"00", (0 + 7722) => x"00", (0 + 7723) => x"00", (0 + 7724) => x"00", (0 + 7725) => x"00", (0 + 7726) => x"00", (0 + 7727) => x"00", (0 + 7728) => x"00", (0 + 7729) => x"00", (0 + 7730) => x"00", (0 + 7731) => x"00", (0 + 7732) => x"00", (0 + 7733) => x"00", (0 + 7734) => x"00", (0 + 7735) => x"00", (0 + 7736) => x"00", (0 + 7737) => x"00", (0 + 7738) => x"00", (0 + 7739) => x"00", (0 + 7740) => x"00", (0 + 7741) => x"00", (0 + 7742) => x"00", (0 + 7743) => x"00", (0 + 7744) => x"00", (0 + 7745) => x"00", (0 + 7746) => x"00", (0 + 7747) => x"00", (0 + 7748) => x"00", (0 + 7749) => x"00", (0 + 7750) => x"00", (0 + 7751) => x"00", (0 + 7752) => x"00", (0 + 7753) => x"00", (0 + 7754) => x"00", (0 + 7755) => x"00", (0 + 7756) => x"00", (0 + 7757) => x"00", (0 + 7758) => x"00", (0 + 7759) => x"00", (0 + 7760) => x"00", (0 + 7761) => x"00", (0 + 7762) => x"00", (0 + 7763) => x"00", (0 + 7764) => x"00", (0 + 7765) => x"00", (0 + 7766) => x"00", (0 + 7767) => x"00", (0 + 7768) => x"00", (0 + 7769) => x"00", (0 + 7770) => x"00", (0 + 7771) => x"00", (0 + 7772) => x"00", (0 + 7773) => x"00", (0 + 7774) => x"00", (0 + 7775) => x"00", (0 + 7776) => x"00", (0 + 7777) => x"00", (0 + 7778) => x"00", (0 + 7779) => x"00", (0 + 7780) => x"00", (0 + 7781) => x"00", (0 + 7782) => x"00", (0 + 7783) => x"00", (0 + 7784) => x"00", (0 + 7785) => x"00", (0 + 7786) => x"00", (0 + 7787) => x"00", (0 + 7788) => x"00", (0 + 7789) => x"00", (0 + 7790) => x"00", (0 + 7791) => x"00", (0 + 7792) => x"00", (0 + 7793) => x"00", (0 + 7794) => x"00", (0 + 7795) => x"00", (0 + 7796) => x"00", (0 + 7797) => x"00", (0 + 7798) => x"00", (0 + 7799) => x"00", (0 + 7800) => x"00", (0 + 7801) => x"00", (0 + 7802) => x"00", (0 + 7803) => x"00", (0 + 7804) => x"00", (0 + 7805) => x"00", (0 + 7806) => x"00", (0 + 7807) => x"00", (0 + 7808) => x"00", (0 + 7809) => x"00", (0 + 7810) => x"00", (0 + 7811) => x"00", (0 + 7812) => x"00", (0 + 7813) => x"00", (0 + 7814) => x"00", (0 + 7815) => x"00", (0 + 7816) => x"00", (0 + 7817) => x"00", (0 + 7818) => x"00", (0 + 7819) => x"00", (0 + 7820) => x"00", (0 + 7821) => x"00", (0 + 7822) => x"00", (0 + 7823) => x"00", (0 + 7824) => x"00", (0 + 7825) => x"00", (0 + 7826) => x"00", (0 + 7827) => x"00", (0 + 7828) => x"00", (0 + 7829) => x"00", (0 + 7830) => x"00", (0 + 7831) => x"00", (0 + 7832) => x"00", (0 + 7833) => x"00", (0 + 7834) => x"00", (0 + 7835) => x"00", (0 + 7836) => x"00", (0 + 7837) => x"00", (0 + 7838) => x"00", (0 + 7839) => x"00", (0 + 7840) => x"00", (0 + 7841) => x"00", (0 + 7842) => x"00", (0 + 7843) => x"00", (0 + 7844) => x"00", (0 + 7845) => x"00", (0 + 7846) => x"00", (0 + 7847) => x"00", (0 + 7848) => x"00", (0 + 7849) => x"00", (0 + 7850) => x"00", (0 + 7851) => x"00", (0 + 7852) => x"00", (0 + 7853) => x"00", (0 + 7854) => x"00", (0 + 7855) => x"00", (0 + 7856) => x"00", (0 + 7857) => x"00", (0 + 7858) => x"00", (0 + 7859) => x"00", (0 + 7860) => x"00", (0 + 7861) => x"00", (0 + 7862) => x"00", (0 + 7863) => x"00", (0 + 7864) => x"00", (0 + 7865) => x"00", (0 + 7866) => x"00", (0 + 7867) => x"00", (0 + 7868) => x"00", (0 + 7869) => x"00", (0 + 7870) => x"00", (0 + 7871) => x"00", (0 + 7872) => x"00", (0 + 7873) => x"00", (0 + 7874) => x"00", (0 + 7875) => x"00", (0 + 7876) => x"00", (0 + 7877) => x"00", (0 + 7878) => x"00", (0 + 7879) => x"00", (0 + 7880) => x"00", (0 + 7881) => x"00", (0 + 7882) => x"00", (0 + 7883) => x"00", (0 + 7884) => x"00", (0 + 7885) => x"00", (0 + 7886) => x"00", (0 + 7887) => x"00", (0 + 7888) => x"00", (0 + 7889) => x"00", (0 + 7890) => x"00", (0 + 7891) => x"00", (0 + 7892) => x"00", (0 + 7893) => x"00", (0 + 7894) => x"00", (0 + 7895) => x"00", (0 + 7896) => x"00", (0 + 7897) => x"00", (0 + 7898) => x"00", (0 + 7899) => x"00", (0 + 7900) => x"00", (0 + 7901) => x"00", (0 + 7902) => x"00", (0 + 7903) => x"00", (0 + 7904) => x"00", (0 + 7905) => x"00", (0 + 7906) => x"00", (0 + 7907) => x"00", (0 + 7908) => x"00", (0 + 7909) => x"00", (0 + 7910) => x"00", (0 + 7911) => x"00", (0 + 7912) => x"00", (0 + 7913) => x"00", (0 + 7914) => x"00", (0 + 7915) => x"00", (0 + 7916) => x"00", (0 + 7917) => x"00", (0 + 7918) => x"00", (0 + 7919) => x"00", (0 + 7920) => x"00", (0 + 7921) => x"00", (0 + 7922) => x"00", (0 + 7923) => x"00", (0 + 7924) => x"00", (0 + 7925) => x"00", (0 + 7926) => x"00", (0 + 7927) => x"00", (0 + 7928) => x"00", (0 + 7929) => x"00", (0 + 7930) => x"00", (0 + 7931) => x"00", (0 + 7932) => x"00", (0 + 7933) => x"00", (0 + 7934) => x"00", (0 + 7935) => x"00", (0 + 7936) => x"00", (0 + 7937) => x"00", (0 + 7938) => x"00", (0 + 7939) => x"00", (0 + 7940) => x"00", (0 + 7941) => x"00", (0 + 7942) => x"00", (0 + 7943) => x"00", (0 + 7944) => x"00", (0 + 7945) => x"00", (0 + 7946) => x"00", (0 + 7947) => x"00", (0 + 7948) => x"00", (0 + 7949) => x"00", (0 + 7950) => x"00", (0 + 7951) => x"00", (0 + 7952) => x"00", (0 + 7953) => x"00", (0 + 7954) => x"00", (0 + 7955) => x"00", (0 + 7956) => x"00", (0 + 7957) => x"00", (0 + 7958) => x"00", (0 + 7959) => x"00", (0 + 7960) => x"00", (0 + 7961) => x"00", (0 + 7962) => x"00", (0 + 7963) => x"00", (0 + 7964) => x"00", (0 + 7965) => x"00", (0 + 7966) => x"00", (0 + 7967) => x"00", (0 + 7968) => x"00", (0 + 7969) => x"00", (0 + 7970) => x"00", (0 + 7971) => x"00", (0 + 7972) => x"00", (0 + 7973) => x"00", (0 + 7974) => x"00", (0 + 7975) => x"00", (0 + 7976) => x"00", (0 + 7977) => x"00", (0 + 7978) => x"00", (0 + 7979) => x"00", (0 + 7980) => x"00", (0 + 7981) => x"00", (0 + 7982) => x"00", (0 + 7983) => x"00", (0 + 7984) => x"00", (0 + 7985) => x"00", (0 + 7986) => x"00", (0 + 7987) => x"00", (0 + 7988) => x"00", (0 + 7989) => x"00", (0 + 7990) => x"00", (0 + 7991) => x"00", (0 + 7992) => x"00", (0 + 7993) => x"00", (0 + 7994) => x"00", (0 + 7995) => x"00", (0 + 7996) => x"00", (0 + 7997) => x"00", (0 + 7998) => x"00", (0 + 7999) => x"00", (0 + 8000) => x"00", (0 + 8001) => x"00", (0 + 8002) => x"00", (0 + 8003) => x"00", (0 + 8004) => x"00", (0 + 8005) => x"00", (0 + 8006) => x"00", (0 + 8007) => x"00", (0 + 8008) => x"00", (0 + 8009) => x"00", (0 + 8010) => x"00", (0 + 8011) => x"00", (0 + 8012) => x"00", (0 + 8013) => x"00", (0 + 8014) => x"00", (0 + 8015) => x"00", (0 + 8016) => x"00", (0 + 8017) => x"00", (0 + 8018) => x"00", (0 + 8019) => x"00", (0 + 8020) => x"00", (0 + 8021) => x"00", (0 + 8022) => x"00", (0 + 8023) => x"00", (0 + 8024) => x"00", (0 + 8025) => x"00", (0 + 8026) => x"00", (0 + 8027) => x"00", (0 + 8028) => x"00", (0 + 8029) => x"00", (0 + 8030) => x"00", (0 + 8031) => x"00", (0 + 8032) => x"00", (0 + 8033) => x"00", (0 + 8034) => x"00", (0 + 8035) => x"00", (0 + 8036) => x"00", (0 + 8037) => x"00", (0 + 8038) => x"00", (0 + 8039) => x"00", (0 + 8040) => x"00", (0 + 8041) => x"00", (0 + 8042) => x"00", (0 + 8043) => x"00", (0 + 8044) => x"00", (0 + 8045) => x"00", (0 + 8046) => x"00", (0 + 8047) => x"00", (0 + 8048) => x"00", (0 + 8049) => x"00", (0 + 8050) => x"00", (0 + 8051) => x"00", (0 + 8052) => x"00", (0 + 8053) => x"00", (0 + 8054) => x"00", (0 + 8055) => x"00", (0 + 8056) => x"00", (0 + 8057) => x"00", (0 + 8058) => x"00", (0 + 8059) => x"00", (0 + 8060) => x"00", (0 + 8061) => x"00", (0 + 8062) => x"00", (0 + 8063) => x"00", (0 + 8064) => x"00", (0 + 8065) => x"00", (0 + 8066) => x"00", (0 + 8067) => x"00", (0 + 8068) => x"00", (0 + 8069) => x"00", (0 + 8070) => x"00", (0 + 8071) => x"00", (0 + 8072) => x"00", (0 + 8073) => x"00", (0 + 8074) => x"00", (0 + 8075) => x"00", (0 + 8076) => x"00", (0 + 8077) => x"00", (0 + 8078) => x"00", (0 + 8079) => x"00", (0 + 8080) => x"00", (0 + 8081) => x"00", (0 + 8082) => x"00", (0 + 8083) => x"00", (0 + 8084) => x"00", (0 + 8085) => x"00", (0 + 8086) => x"00", (0 + 8087) => x"00", (0 + 8088) => x"00", (0 + 8089) => x"00", (0 + 8090) => x"00", (0 + 8091) => x"00", (0 + 8092) => x"00", (0 + 8093) => x"00", (0 + 8094) => x"00", (0 + 8095) => x"00", (0 + 8096) => x"00", (0 + 8097) => x"00", (0 + 8098) => x"00", (0 + 8099) => x"00", (0 + 8100) => x"00", (0 + 8101) => x"00", (0 + 8102) => x"00", (0 + 8103) => x"00", (0 + 8104) => x"00", (0 + 8105) => x"00", (0 + 8106) => x"00", (0 + 8107) => x"00", (0 + 8108) => x"00", (0 + 8109) => x"00", (0 + 8110) => x"00", (0 + 8111) => x"00", (0 + 8112) => x"00", (0 + 8113) => x"00", (0 + 8114) => x"00", (0 + 8115) => x"00", (0 + 8116) => x"00", (0 + 8117) => x"00", (0 + 8118) => x"00", (0 + 8119) => x"00", (0 + 8120) => x"00", (0 + 8121) => x"00", (0 + 8122) => x"00", (0 + 8123) => x"00", (0 + 8124) => x"00", (0 + 8125) => x"00", (0 + 8126) => x"00", (0 + 8127) => x"00", (0 + 8128) => x"00", (0 + 8129) => x"00", (0 + 8130) => x"00", (0 + 8131) => x"00", (0 + 8132) => x"00", (0 + 8133) => x"00", (0 + 8134) => x"00", (0 + 8135) => x"00", (0 + 8136) => x"00", (0 + 8137) => x"00", (0 + 8138) => x"00", (0 + 8139) => x"00", (0 + 8140) => x"00", (0 + 8141) => x"00", (0 + 8142) => x"00", (0 + 8143) => x"00", (0 + 8144) => x"00", (0 + 8145) => x"00", (0 + 8146) => x"00", (0 + 8147) => x"00", (0 + 8148) => x"00", (0 + 8149) => x"00", (0 + 8150) => x"00", (0 + 8151) => x"00", (0 + 8152) => x"00", (0 + 8153) => x"00", (0 + 8154) => x"00", (0 + 8155) => x"00", (0 + 8156) => x"00", (0 + 8157) => x"00", (0 + 8158) => x"00", (0 + 8159) => x"00", (0 + 8160) => x"00", (0 + 8161) => x"00", (0 + 8162) => x"00", (0 + 8163) => x"00", (0 + 8164) => x"00", (0 + 8165) => x"00", (0 + 8166) => x"00", (0 + 8167) => x"00", (0 + 8168) => x"00", (0 + 8169) => x"00", (0 + 8170) => x"00", (0 + 8171) => x"00", (0 + 8172) => x"00", (0 + 8173) => x"00", (0 + 8174) => x"00", (0 + 8175) => x"00", (0 + 8176) => x"00", (0 + 8177) => x"00", (0 + 8178) => x"00", (0 + 8179) => x"00", (0 + 8180) => x"00", (0 + 8181) => x"00", (0 + 8182) => x"00", (0 + 8183) => x"00", (0 + 8184) => x"00", (0 + 8185) => x"00", (0 + 8186) => x"00", (0 + 8187) => x"00", (0 + 8188) => x"00", (0 + 8189) => x"00", (0 + 8190) => x"00", (0 + 8191) => x"00", 