library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity stub_ram_0 is
    Port ( 
           address : in STD_LOGIC_VECTOR (11 downto 0);
           clock : in STD_LOGIC;
           we : in STD_LOGIC;
           dataIn : in STD_LOGIC_VECTOR (7 downto 0);
           dataOut : out STD_LOGIC_VECTOR (7 downto 0));
end stub_ram_0;

architecture Behavioral of stub_ram_0 is
    type RAM is array ( ( 4 * 1024 ) - 1 downto 0 ) of std_logic_vector( 7 downto 0 );
    
    signal sys_RAM : RAM := (
                                (0 + 0) => x"37", (0 + 1) => x"6f", (0 + 2) => x"13", (0 + 3) => x"93", (0 + 4) => x"37", (0 + 5) => x"23", (0 + 6) => x"23", (0 + 7) => x"23", (0 + 8) => x"23", (0 + 9) => x"33", (0 + 10) => x"23", (0 + 11) => x"23", (0 + 12) => x"23", (0 + 13) => x"b7", (0 + 14) => x"23", (0 + 15) => x"97", (0 + 16) => x"93", (0 + 17) => x"17", (0 + 18) => x"13", (0 + 19) => x"13", (0 + 20) => x"93", (0 + 21) => x"13", (0 + 22) => x"13", (0 + 23) => x"93", (0 + 24) => x"93", (0 + 25) => x"13", (0 + 26) => x"93", (0 + 27) => x"37", (0 + 28) => x"93", (0 + 29) => x"b7", (0 + 30) => x"93", (0 + 31) => x"13", (0 + 32) => x"93", (0 + 33) => x"97", (0 + 34) => x"23", (0 + 35) => x"97", (0 + 36) => x"23", (0 + 37) => x"03", (0 + 38) => x"97", (0 + 39) => x"93", (0 + 40) => x"33", (0 + 41) => x"23", (0 + 42) => x"93", (0 + 43) => x"03", (0 + 44) => x"e3", (0 + 45) => x"03", (0 + 46) => x"b3", (0 + 47) => x"83", (0 + 48) => x"13", (0 + 49) => x"63", (0 + 50) => x"13", (0 + 51) => x"83", (0 + 52) => x"e3", (0 + 53) => x"33", (0 + 54) => x"93", (0 + 55) => x"b3", (0 + 56) => x"13", (0 + 57) => x"63", (0 + 58) => x"97", (0 + 59) => x"23", (0 + 60) => x"13", (0 + 61) => x"e3", (0 + 62) => x"97", (0 + 63) => x"23", (0 + 64) => x"97", (0 + 65) => x"23", (0 + 66) => x"97", (0 + 67) => x"23", (0 + 68) => x"93", (0 + 69) => x"b3", (0 + 70) => x"23", (0 + 71) => x"93", (0 + 72) => x"e3", (0 + 73) => x"97", (0 + 74) => x"93", (0 + 75) => x"93", (0 + 76) => x"03", (0 + 77) => x"e3", (0 + 78) => x"b3", (0 + 79) => x"13", (0 + 80) => x"93", (0 + 81) => x"63", (0 + 82) => x"17", (0 + 83) => x"23", (0 + 84) => x"93", (0 + 85) => x"e3", (0 + 86) => x"97", (0 + 87) => x"93", (0 + 88) => x"93", (0 + 89) => x"03", (0 + 90) => x"e3", (0 + 91) => x"b3", (0 + 92) => x"b3", (0 + 93) => x"13", (0 + 94) => x"63", (0 + 95) => x"97", (0 + 96) => x"23", (0 + 97) => x"13", (0 + 98) => x"e3", (0 + 99) => x"97", (0 + 100) => x"23", (0 + 101) => x"97", (0 + 102) => x"93", (0 + 103) => x"93", (0 + 104) => x"03", (0 + 105) => x"e3", (0 + 106) => x"33", (0 + 107) => x"b3", (0 + 108) => x"b3", (0 + 109) => x"13", (0 + 110) => x"63", (0 + 111) => x"97", (0 + 112) => x"23", (0 + 113) => x"13", (0 + 114) => x"e3", (0 + 115) => x"23", (0 + 116) => x"23", (0 + 117) => x"83", (0 + 118) => x"23", (0 + 119) => x"93", (0 + 120) => x"93", (0 + 121) => x"13", (0 + 122) => x"63", (0 + 123) => x"93", (0 + 124) => x"b3", (0 + 125) => x"b3", (0 + 126) => x"6f", (0 + 127) => x"13", (0 + 128) => x"63", (0 + 129) => x"93", (0 + 130) => x"b3", (0 + 131) => x"b3", (0 + 132) => x"6f", (0 + 133) => x"13", (0 + 134) => x"63", (0 + 135) => x"13", (0 + 136) => x"13", (0 + 137) => x"e3", (0 + 138) => x"13", (0 + 139) => x"13", (0 + 140) => x"6f", (0 + 141) => x"13", (0 + 142) => x"6f", (0 + 143) => x"13", (0 + 144) => x"63", (0 + 145) => x"13", (0 + 146) => x"13", (0 + 147) => x"e3", (0 + 148) => x"13", (0 + 149) => x"13", (0 + 150) => x"6f", (0 + 151) => x"93", (0 + 152) => x"63", (0 + 153) => x"83", (0 + 154) => x"23", (0 + 155) => x"03", (0 + 156) => x"83", (0 + 157) => x"03", (0 + 158) => x"83", (0 + 159) => x"03", (0 + 160) => x"83", (0 + 161) => x"03", (0 + 162) => x"13", (0 + 163) => x"67", (0 + 164) => x"b7", (0 + 165) => x"23", (0 + 166) => x"93", (0 + 167) => x"97", (0 + 168) => x"23", (0 + 169) => x"97", (0 + 170) => x"23", (0 + 171) => x"03", (0 + 172) => x"17", (0 + 173) => x"13", (0 + 174) => x"13", (0 + 175) => x"33", (0 + 176) => x"93", (0 + 177) => x"23", (0 + 178) => x"93", (0 + 179) => x"03", (0 + 180) => x"e3", (0 + 181) => x"03", (0 + 182) => x"b3", (0 + 183) => x"83", (0 + 184) => x"13", (0 + 185) => x"63", (0 + 186) => x"13", (0 + 187) => x"83", (0 + 188) => x"e3", (0 + 189) => x"33", (0 + 190) => x"93", (0 + 191) => x"b3", (0 + 192) => x"93", (0 + 193) => x"13", (0 + 194) => x"63", (0 + 195) => x"93", (0 + 196) => x"93", (0 + 197) => x"17", (0 + 198) => x"23", (0 + 199) => x"13", (0 + 200) => x"e3", (0 + 201) => x"93", (0 + 202) => x"17", (0 + 203) => x"23", (0 + 204) => x"17", (0 + 205) => x"23", (0 + 206) => x"b7", (0 + 207) => x"13", (0 + 208) => x"33", (0 + 209) => x"17", (0 + 210) => x"23", (0 + 211) => x"93", (0 + 212) => x"b3", (0 + 213) => x"13", (0 + 214) => x"93", (0 + 215) => x"23", (0 + 216) => x"93", (0 + 217) => x"e3", (0 + 218) => x"97", (0 + 219) => x"93", (0 + 220) => x"93", (0 + 221) => x"93", (0 + 222) => x"03", (0 + 223) => x"e3", (0 + 224) => x"b3", (0 + 225) => x"93", (0 + 226) => x"13", (0 + 227) => x"93", (0 + 228) => x"63", (0 + 229) => x"93", (0 + 230) => x"13", (0 + 231) => x"17", (0 + 232) => x"23", (0 + 233) => x"93", (0 + 234) => x"e3", (0 + 235) => x"93", (0 + 236) => x"17", (0 + 237) => x"23", (0 + 238) => x"13", (0 + 239) => x"b7", (0 + 240) => x"23", (0 + 241) => x"23", (0 + 242) => x"b7", (0 + 243) => x"23", (0 + 244) => x"13", (0 + 245) => x"67", (0 + 246) => x"13", (0 + 247) => x"6f", (0 + 248) => x"17", (0 + 249) => x"23", (0 + 250) => x"37", (0 + 251) => x"13", (0 + 252) => x"97", (0 + 253) => x"93", (0 + 254) => x"13", (0 + 255) => x"97", (0 + 256) => x"23", (0 + 257) => x"23", (0 + 258) => x"23", (0 + 259) => x"23", (0 + 260) => x"97", (0 + 261) => x"93", (0 + 262) => x"23", (0 + 263) => x"23", (0 + 264) => x"23", (0 + 265) => x"23", (0 + 266) => x"23", (0 + 267) => x"23", (0 + 268) => x"23", (0 + 269) => x"23", (0 + 270) => x"23", (0 + 271) => x"23", (0 + 272) => x"23", (0 + 273) => x"23", (0 + 274) => x"13", (0 + 275) => x"13", (0 + 276) => x"93", (0 + 277) => x"93", (0 + 278) => x"93", (0 + 279) => x"b3", (0 + 280) => x"23", (0 + 281) => x"a3", (0 + 282) => x"93", (0 + 283) => x"23", (0 + 284) => x"13", (0 + 285) => x"13", (0 + 286) => x"a3", (0 + 287) => x"13", (0 + 288) => x"13", (0 + 289) => x"13", (0 + 290) => x"13", (0 + 291) => x"63", (0 + 292) => x"23", (0 + 293) => x"63", (0 + 294) => x"a3", (0 + 295) => x"63", (0 + 296) => x"23", (0 + 297) => x"63", (0 + 298) => x"a3", (0 + 299) => x"13", (0 + 300) => x"e3", (0 + 301) => x"23", (0 + 302) => x"a3", (0 + 303) => x"23", (0 + 304) => x"a3", (0 + 305) => x"b7", (0 + 306) => x"23", (0 + 307) => x"b7", (0 + 308) => x"37", (0 + 309) => x"93", (0 + 310) => x"23", (0 + 311) => x"13", (0 + 312) => x"b7", (0 + 313) => x"23", (0 + 314) => x"13", (0 + 315) => x"13", (0 + 316) => x"93", (0 + 317) => x"13", (0 + 318) => x"13", (0 + 319) => x"93", (0 + 320) => x"b7", (0 + 321) => x"b7", (0 + 322) => x"13", (0 + 323) => x"13", (0 + 324) => x"b7", (0 + 325) => x"13", (0 + 326) => x"b3", (0 + 327) => x"93", (0 + 328) => x"23", (0 + 329) => x"33", (0 + 330) => x"93", (0 + 331) => x"b3", (0 + 332) => x"83", (0 + 333) => x"13", (0 + 334) => x"b3", (0 + 335) => x"93", (0 + 336) => x"13", (0 + 337) => x"b3", (0 + 338) => x"33", (0 + 339) => x"23", (0 + 340) => x"b3", (0 + 341) => x"93", (0 + 342) => x"83", (0 + 343) => x"13", (0 + 344) => x"23", (0 + 345) => x"b3", (0 + 346) => x"83", (0 + 347) => x"17", (0 + 348) => x"23", (0 + 349) => x"97", (0 + 350) => x"23", (0 + 351) => x"13", (0 + 352) => x"93", (0 + 353) => x"33", (0 + 354) => x"b3", (0 + 355) => x"97", (0 + 356) => x"23", (0 + 357) => x"23", (0 + 358) => x"b3", (0 + 359) => x"93", (0 + 360) => x"23", (0 + 361) => x"b3", (0 + 362) => x"03", (0 + 363) => x"97", (0 + 364) => x"23", (0 + 365) => x"93", (0 + 366) => x"b3", (0 + 367) => x"93", (0 + 368) => x"33", (0 + 369) => x"b3", (0 + 370) => x"93", (0 + 371) => x"23", (0 + 372) => x"b3", (0 + 373) => x"13", (0 + 374) => x"13", (0 + 375) => x"93", (0 + 376) => x"b3", (0 + 377) => x"23", (0 + 378) => x"93", (0 + 379) => x"13", (0 + 380) => x"93", (0 + 381) => x"93", (0 + 382) => x"b3", (0 + 383) => x"b3", (0 + 384) => x"33", (0 + 385) => x"b3", (0 + 386) => x"13", (0 + 387) => x"13", (0 + 388) => x"b3", (0 + 389) => x"33", (0 + 390) => x"b3", (0 + 391) => x"b3", (0 + 392) => x"63", (0 + 393) => x"13", (0 + 394) => x"23", (0 + 395) => x"33", (0 + 396) => x"33", (0 + 397) => x"b3", (0 + 398) => x"e3", (0 + 399) => x"97", (0 + 400) => x"93", (0 + 401) => x"13", (0 + 402) => x"b7", (0 + 403) => x"13", (0 + 404) => x"93", (0 + 405) => x"93", (0 + 406) => x"23", (0 + 407) => x"13", (0 + 408) => x"93", (0 + 409) => x"13", (0 + 410) => x"13", (0 + 411) => x"97", (0 + 412) => x"23", (0 + 413) => x"97", (0 + 414) => x"23", (0 + 415) => x"97", (0 + 416) => x"93", (0 + 417) => x"93", (0 + 418) => x"03", (0 + 419) => x"e3", (0 + 420) => x"b3", (0 + 421) => x"13", (0 + 422) => x"93", (0 + 423) => x"63", (0 + 424) => x"17", (0 + 425) => x"23", (0 + 426) => x"93", (0 + 427) => x"e3", (0 + 428) => x"63", (0 + 429) => x"13", (0 + 430) => x"33", (0 + 431) => x"13", (0 + 432) => x"33", (0 + 433) => x"13", (0 + 434) => x"13", (0 + 435) => x"63", (0 + 436) => x"97", (0 + 437) => x"23", (0 + 438) => x"13", (0 + 439) => x"13", (0 + 440) => x"e3", (0 + 441) => x"b7", (0 + 442) => x"13", (0 + 443) => x"23", (0 + 444) => x"23", (0 + 445) => x"83", (0 + 446) => x"37", (0 + 447) => x"23", (0 + 448) => x"93", (0 + 449) => x"93", (0 + 450) => x"13", (0 + 451) => x"63", (0 + 452) => x"93", (0 + 453) => x"e3", (0 + 454) => x"13", (0 + 455) => x"e3", (0 + 456) => x"93", (0 + 457) => x"13", (0 + 458) => x"6f", (0 + 459) => x"63", (0 + 460) => x"97", (0 + 461) => x"23", (0 + 462) => x"83", (0 + 463) => x"b3", (0 + 464) => x"23", (0 + 465) => x"83", (0 + 466) => x"83", (0 + 467) => x"63", (0 + 468) => x"93", (0 + 469) => x"93", (0 + 470) => x"83", (0 + 471) => x"e3", (0 + 472) => x"b3", (0 + 473) => x"93", (0 + 474) => x"93", (0 + 475) => x"63", (0 + 476) => x"6f", (0 + 477) => x"93", (0 + 478) => x"97", (0 + 479) => x"23", (0 + 480) => x"93", (0 + 481) => x"e3", (0 + 482) => x"6f", (0 + 483) => x"13", (0 + 484) => x"63", (0 + 485) => x"e3", (0 + 486) => x"13", (0 + 487) => x"e3", (0 + 488) => x"93", (0 + 489) => x"13", (0 + 490) => x"6f", (0 + 491) => x"93", (0 + 492) => x"6f", (0 + 493) => x"93", (0 + 494) => x"e3", (0 + 495) => x"93", (0 + 496) => x"b3", (0 + 497) => x"93", (0 + 498) => x"b3", (0 + 499) => x"03", (0 + 500) => x"03", (0 + 501) => x"e7", (0 + 502) => x"6f", (0 + 503) => x"97", (0 + 504) => x"23", (0 + 505) => x"6f", (0 + 506) => x"00", (0 + 507) => x"c8", (0 + 508) => x"90", (0 + 509) => x"44", (0 + 510) => x"dc", (0 + 511) => x"90", (0 + 512) => x"4c", (0 + 513) => x"f0", (0 + 514) => x"08", (0 + 515) => x"4c", (0 + 516) => x"04", (0 + 517) => x"90", (0 + 518) => x"54", (0 + 519) => x"18", (0 + 520) => x"08", (0 + 521) => x"54", (0 + 522) => x"30", (0 + 523) => x"34", (0 + 524) => x"38", (0 + 525) => x"43", (0 + 526) => x"98", (0 + 527) => x"ec", (0 + 528) => x"05", (0 + 529) => x"d0", (0 + 530) => x"2c", (0 + 531) => x"f8", (0 + 532) => x"00", (0 + 533) => x"20", (0 + 534) => x"04", (0 + 535) => x"53", (0 + 536) => x"20", (0 + 537) => x"56", (0 + 538) => x"45", (0 + 539) => x"20", (0 + 540) => x"20", (0 + 541) => x"20", (0 + 542) => x"20", (0 + 543) => x"20", (0 + 544) => x"20", (0 + 545) => x"00", (0 + 546) => x"58", (0 + 547) => x"20", (0 + 548) => x"4e", (0 + 549) => x"20", (0 + 550) => x"4d", (0 + 551) => x"20", (0 + 552) => x"55", (0 + 553) => x"53", (0 + 554) => x"54", (0 + 555) => x"20", (0 + 556) => x"20", (0 + 557) => x"20", (0 + 558) => x"20", (0 + 559) => x"20", (0 + 560) => x"20", (0 + 561) => x"20", (0 + 562) => x"31", (0 + 563) => x"68", (0 + 564) => x"6d", (0 + 565) => x"61", (0 + 566) => x"6f", (0 + 567) => x"32", (0 + 568) => x"68", (0 + 569) => x"6d", (0 + 570) => x"61", (0 + 571) => x"61", (0 + 572) => x"33", (0 + 573) => x"65", (0 + 574) => x"6d", (0 + 575) => x"61", (0 + 576) => x"61", (0 + 577) => x"34", (0 + 578) => x"68", (0 + 579) => x"6d", (0 + 580) => x"61", (0 + 581) => x"61", (0 + 582) => x"35", (0 + 583) => x"65", (0 + 584) => x"6d", (0 + 585) => x"61", (0 + 586) => x"61", (0 + 587) => x"ef", (0 + 588) => x"00", (0 + 589) => x"00", (0 + 590) => x"00", (0 + 591) => x"00", (0 + 592) => x"00", (0 + 593) => x"00", (0 + 594) => x"00", (0 + 595) => x"00", (0 + 596) => x"00", (0 + 597) => x"00", (0 + 598) => x"00", (0 + 599) => x"00", (0 + 600) => x"00", (0 + 601) => x"00", (0 + 602) => x"00", (0 + 603) => x"00", (0 + 604) => x"00", (0 + 605) => x"00", (0 + 606) => x"00", (0 + 607) => x"00", (0 + 608) => x"00", (0 + 609) => x"00", (0 + 610) => x"00", (0 + 611) => x"00", (0 + 612) => x"00", (0 + 613) => x"00", (0 + 614) => x"00", (0 + 615) => x"00", (0 + 616) => x"00", (0 + 617) => x"00", (0 + 618) => x"00", (0 + 619) => x"00", (0 + 620) => x"00", (0 + 621) => x"00", (0 + 622) => x"00", (0 + 623) => x"00", (0 + 624) => x"00", (0 + 625) => x"00", (0 + 626) => x"00", (0 + 627) => x"00", (0 + 628) => x"00", (0 + 629) => x"00", (0 + 630) => x"00", (0 + 631) => x"00", (0 + 632) => x"00", (0 + 633) => x"00", (0 + 634) => x"00", (0 + 635) => x"00", (0 + 636) => x"00", (0 + 637) => x"00", (0 + 638) => x"00", (0 + 639) => x"00", (0 + 640) => x"00", (0 + 641) => x"00", (0 + 642) => x"00", (0 + 643) => x"00", (0 + 644) => x"00", (0 + 645) => x"00", (0 + 646) => x"00", (0 + 647) => x"00", (0 + 648) => x"00", (0 + 649) => x"00", (0 + 650) => x"00", (0 + 651) => x"00", (0 + 652) => x"00", (0 + 653) => x"00", (0 + 654) => x"00", (0 + 655) => x"00", (0 + 656) => x"00", (0 + 657) => x"00", (0 + 658) => x"00", (0 + 659) => x"00", (0 + 660) => x"00", (0 + 661) => x"00", (0 + 662) => x"00", (0 + 663) => x"00", (0 + 664) => x"00", (0 + 665) => x"00", (0 + 666) => x"00", (0 + 667) => x"00", (0 + 668) => x"00", (0 + 669) => x"00", (0 + 670) => x"00", (0 + 671) => x"00", (0 + 672) => x"00", (0 + 673) => x"00", (0 + 674) => x"00", (0 + 675) => x"00", (0 + 676) => x"00", (0 + 677) => x"00", (0 + 678) => x"00", (0 + 679) => x"00", (0 + 680) => x"00", (0 + 681) => x"00", (0 + 682) => x"00", (0 + 683) => x"00", (0 + 684) => x"00", (0 + 685) => x"00", (0 + 686) => x"00", (0 + 687) => x"00", (0 + 688) => x"00", (0 + 689) => x"00", (0 + 690) => x"00", (0 + 691) => x"00", (0 + 692) => x"00", (0 + 693) => x"00", (0 + 694) => x"00", (0 + 695) => x"00", (0 + 696) => x"00", (0 + 697) => x"00", (0 + 698) => x"00", (0 + 699) => x"00", (0 + 700) => x"00", (0 + 701) => x"00", (0 + 702) => x"00", (0 + 703) => x"00", (0 + 704) => x"00", (0 + 705) => x"00", (0 + 706) => x"00", (0 + 707) => x"00", (0 + 708) => x"00", (0 + 709) => x"00", (0 + 710) => x"00", (0 + 711) => x"00", (0 + 712) => x"00", (0 + 713) => x"00", (0 + 714) => x"00", (0 + 715) => x"00", (0 + 716) => x"00", (0 + 717) => x"00", (0 + 718) => x"00", (0 + 719) => x"00", (0 + 720) => x"00", (0 + 721) => x"00", (0 + 722) => x"00", (0 + 723) => x"00", (0 + 724) => x"00", (0 + 725) => x"00", (0 + 726) => x"00", (0 + 727) => x"00", (0 + 728) => x"00", (0 + 729) => x"00", (0 + 730) => x"00", (0 + 731) => x"00", (0 + 732) => x"00", (0 + 733) => x"00", (0 + 734) => x"00", (0 + 735) => x"00", (0 + 736) => x"00", (0 + 737) => x"00", (0 + 738) => x"00", (0 + 739) => x"00", (0 + 740) => x"00", (0 + 741) => x"00", (0 + 742) => x"00", (0 + 743) => x"00", (0 + 744) => x"00", (0 + 745) => x"00", (0 + 746) => x"00", (0 + 747) => x"00", (0 + 748) => x"00", (0 + 749) => x"00", (0 + 750) => x"00", (0 + 751) => x"00", (0 + 752) => x"00", (0 + 753) => x"00", (0 + 754) => x"00", (0 + 755) => x"00", (0 + 756) => x"00", (0 + 757) => x"00", (0 + 758) => x"00", (0 + 759) => x"00", (0 + 760) => x"00", (0 + 761) => x"00", (0 + 762) => x"00", (0 + 763) => x"00", (0 + 764) => x"00", (0 + 765) => x"00", (0 + 766) => x"00", (0 + 767) => x"00", (0 + 768) => x"00", (0 + 769) => x"00", (0 + 770) => x"00", (0 + 771) => x"00", (0 + 772) => x"00", (0 + 773) => x"00", (0 + 774) => x"00", (0 + 775) => x"00", (0 + 776) => x"00", (0 + 777) => x"00", (0 + 778) => x"00", (0 + 779) => x"00", (0 + 780) => x"00", (0 + 781) => x"00", (0 + 782) => x"00", (0 + 783) => x"00", (0 + 784) => x"00", (0 + 785) => x"00", (0 + 786) => x"00", (0 + 787) => x"00", (0 + 788) => x"00", (0 + 789) => x"00", (0 + 790) => x"00", (0 + 791) => x"00", (0 + 792) => x"00", (0 + 793) => x"00", (0 + 794) => x"00", (0 + 795) => x"00", (0 + 796) => x"00", (0 + 797) => x"00", (0 + 798) => x"00", (0 + 799) => x"00", (0 + 800) => x"00", (0 + 801) => x"00", (0 + 802) => x"00", (0 + 803) => x"00", (0 + 804) => x"00", (0 + 805) => x"00", (0 + 806) => x"00", (0 + 807) => x"00", (0 + 808) => x"00", (0 + 809) => x"00", (0 + 810) => x"00", (0 + 811) => x"00", (0 + 812) => x"00", (0 + 813) => x"00", (0 + 814) => x"00", (0 + 815) => x"00", (0 + 816) => x"00", (0 + 817) => x"00", (0 + 818) => x"00", (0 + 819) => x"00", (0 + 820) => x"00", (0 + 821) => x"00", (0 + 822) => x"00", (0 + 823) => x"00", (0 + 824) => x"00", (0 + 825) => x"00", (0 + 826) => x"00", (0 + 827) => x"00", (0 + 828) => x"00", (0 + 829) => x"00", (0 + 830) => x"00", (0 + 831) => x"00", (0 + 832) => x"00", (0 + 833) => x"00", (0 + 834) => x"00", (0 + 835) => x"00", (0 + 836) => x"00", (0 + 837) => x"00", (0 + 838) => x"00", (0 + 839) => x"00", (0 + 840) => x"00", (0 + 841) => x"00", (0 + 842) => x"00", (0 + 843) => x"00", (0 + 844) => x"00", (0 + 845) => x"00", (0 + 846) => x"00", (0 + 847) => x"00", (0 + 848) => x"00", (0 + 849) => x"00", (0 + 850) => x"00", (0 + 851) => x"00", (0 + 852) => x"00", (0 + 853) => x"00", (0 + 854) => x"00", (0 + 855) => x"00", (0 + 856) => x"00", (0 + 857) => x"00", (0 + 858) => x"00", (0 + 859) => x"00", (0 + 860) => x"00", (0 + 861) => x"00", (0 + 862) => x"00", (0 + 863) => x"00", (0 + 864) => x"00", (0 + 865) => x"00", (0 + 866) => x"00", (0 + 867) => x"00", (0 + 868) => x"00", (0 + 869) => x"00", (0 + 870) => x"00", (0 + 871) => x"00", (0 + 872) => x"00", (0 + 873) => x"00", (0 + 874) => x"00", (0 + 875) => x"00", (0 + 876) => x"00", (0 + 877) => x"00", (0 + 878) => x"00", (0 + 879) => x"00", (0 + 880) => x"00", (0 + 881) => x"00", (0 + 882) => x"00", (0 + 883) => x"00", (0 + 884) => x"00", (0 + 885) => x"00", (0 + 886) => x"00", (0 + 887) => x"00", (0 + 888) => x"00", (0 + 889) => x"00", (0 + 890) => x"00", (0 + 891) => x"00", (0 + 892) => x"00", (0 + 893) => x"00", (0 + 894) => x"00", (0 + 895) => x"00", (0 + 896) => x"00", (0 + 897) => x"00", (0 + 898) => x"00", (0 + 899) => x"00", (0 + 900) => x"00", (0 + 901) => x"00", (0 + 902) => x"00", (0 + 903) => x"00", (0 + 904) => x"00", (0 + 905) => x"00", (0 + 906) => x"00", (0 + 907) => x"00", (0 + 908) => x"00", (0 + 909) => x"00", (0 + 910) => x"00", (0 + 911) => x"00", (0 + 912) => x"00", (0 + 913) => x"00", (0 + 914) => x"00", (0 + 915) => x"00", (0 + 916) => x"00", (0 + 917) => x"00", (0 + 918) => x"00", (0 + 919) => x"00", (0 + 920) => x"00", (0 + 921) => x"00", (0 + 922) => x"00", (0 + 923) => x"00", (0 + 924) => x"00", (0 + 925) => x"00", (0 + 926) => x"00", (0 + 927) => x"00", (0 + 928) => x"00", (0 + 929) => x"00", (0 + 930) => x"00", (0 + 931) => x"00", (0 + 932) => x"00", (0 + 933) => x"00", (0 + 934) => x"00", (0 + 935) => x"00", (0 + 936) => x"00", (0 + 937) => x"00", (0 + 938) => x"00", (0 + 939) => x"00", (0 + 940) => x"00", (0 + 941) => x"00", (0 + 942) => x"00", (0 + 943) => x"00", (0 + 944) => x"00", (0 + 945) => x"00", (0 + 946) => x"00", (0 + 947) => x"00", (0 + 948) => x"00", (0 + 949) => x"00", (0 + 950) => x"00", (0 + 951) => x"00", (0 + 952) => x"00", (0 + 953) => x"00", (0 + 954) => x"00", (0 + 955) => x"00", (0 + 956) => x"00", (0 + 957) => x"00", (0 + 958) => x"00", (0 + 959) => x"00", (0 + 960) => x"00", (0 + 961) => x"00", (0 + 962) => x"00", (0 + 963) => x"00", (0 + 964) => x"00", (0 + 965) => x"00", (0 + 966) => x"00", (0 + 967) => x"00", (0 + 968) => x"00", (0 + 969) => x"00", (0 + 970) => x"00", (0 + 971) => x"00", (0 + 972) => x"00", (0 + 973) => x"00", (0 + 974) => x"00", (0 + 975) => x"00", (0 + 976) => x"00", (0 + 977) => x"00", (0 + 978) => x"00", (0 + 979) => x"00", (0 + 980) => x"00", (0 + 981) => x"00", (0 + 982) => x"00", (0 + 983) => x"00", (0 + 984) => x"00", (0 + 985) => x"00", (0 + 986) => x"00", (0 + 987) => x"00", (0 + 988) => x"00", (0 + 989) => x"00", (0 + 990) => x"00", (0 + 991) => x"00", (0 + 992) => x"00", (0 + 993) => x"00", (0 + 994) => x"00", (0 + 995) => x"00", (0 + 996) => x"00", (0 + 997) => x"00", (0 + 998) => x"00", (0 + 999) => x"00", (0 + 1000) => x"00", (0 + 1001) => x"00", (0 + 1002) => x"00", (0 + 1003) => x"00", (0 + 1004) => x"00", (0 + 1005) => x"00", (0 + 1006) => x"00", (0 + 1007) => x"00", (0 + 1008) => x"00", (0 + 1009) => x"00", (0 + 1010) => x"00", (0 + 1011) => x"00", (0 + 1012) => x"00", (0 + 1013) => x"00", (0 + 1014) => x"00", (0 + 1015) => x"00", (0 + 1016) => x"00", (0 + 1017) => x"00", (0 + 1018) => x"00", (0 + 1019) => x"00", (0 + 1020) => x"00", (0 + 1021) => x"00", (0 + 1022) => x"00", (0 + 1023) => x"00", (0 + 1024) => x"00", (0 + 1025) => x"00", (0 + 1026) => x"00", (0 + 1027) => x"00", (0 + 1028) => x"00", (0 + 1029) => x"00", (0 + 1030) => x"00", (0 + 1031) => x"00", (0 + 1032) => x"00", (0 + 1033) => x"00", (0 + 1034) => x"00", (0 + 1035) => x"00", (0 + 1036) => x"00", (0 + 1037) => x"00", (0 + 1038) => x"00", (0 + 1039) => x"00", (0 + 1040) => x"00", (0 + 1041) => x"00", (0 + 1042) => x"00", (0 + 1043) => x"00", (0 + 1044) => x"00", (0 + 1045) => x"00", (0 + 1046) => x"00", (0 + 1047) => x"00", (0 + 1048) => x"00", (0 + 1049) => x"00", (0 + 1050) => x"00", (0 + 1051) => x"00", (0 + 1052) => x"00", (0 + 1053) => x"00", (0 + 1054) => x"00", (0 + 1055) => x"00", (0 + 1056) => x"00", (0 + 1057) => x"00", (0 + 1058) => x"00", (0 + 1059) => x"00", (0 + 1060) => x"00", (0 + 1061) => x"00", (0 + 1062) => x"00", (0 + 1063) => x"00", (0 + 1064) => x"00", (0 + 1065) => x"00", (0 + 1066) => x"00", (0 + 1067) => x"00", (0 + 1068) => x"00", (0 + 1069) => x"00", (0 + 1070) => x"00", (0 + 1071) => x"00", (0 + 1072) => x"00", (0 + 1073) => x"00", (0 + 1074) => x"00", (0 + 1075) => x"00", (0 + 1076) => x"00", (0 + 1077) => x"00", (0 + 1078) => x"00", (0 + 1079) => x"00", (0 + 1080) => x"00", (0 + 1081) => x"00", (0 + 1082) => x"00", (0 + 1083) => x"00", (0 + 1084) => x"00", (0 + 1085) => x"00", (0 + 1086) => x"00", (0 + 1087) => x"00", (0 + 1088) => x"00", (0 + 1089) => x"00", (0 + 1090) => x"00", (0 + 1091) => x"00", (0 + 1092) => x"00", (0 + 1093) => x"00", (0 + 1094) => x"00", (0 + 1095) => x"00", (0 + 1096) => x"00", (0 + 1097) => x"00", (0 + 1098) => x"00", (0 + 1099) => x"00", (0 + 1100) => x"00", (0 + 1101) => x"00", (0 + 1102) => x"00", (0 + 1103) => x"00", (0 + 1104) => x"00", (0 + 1105) => x"00", (0 + 1106) => x"00", (0 + 1107) => x"00", (0 + 1108) => x"00", (0 + 1109) => x"00", (0 + 1110) => x"00", (0 + 1111) => x"00", (0 + 1112) => x"00", (0 + 1113) => x"00", (0 + 1114) => x"00", (0 + 1115) => x"00", (0 + 1116) => x"00", (0 + 1117) => x"00", (0 + 1118) => x"00", (0 + 1119) => x"00", (0 + 1120) => x"00", (0 + 1121) => x"00", (0 + 1122) => x"00", (0 + 1123) => x"00", (0 + 1124) => x"00", (0 + 1125) => x"00", (0 + 1126) => x"00", (0 + 1127) => x"00", (0 + 1128) => x"00", (0 + 1129) => x"00", (0 + 1130) => x"00", (0 + 1131) => x"00", (0 + 1132) => x"00", (0 + 1133) => x"00", (0 + 1134) => x"00", (0 + 1135) => x"00", (0 + 1136) => x"00", (0 + 1137) => x"00", (0 + 1138) => x"00", (0 + 1139) => x"00", (0 + 1140) => x"00", (0 + 1141) => x"00", (0 + 1142) => x"00", (0 + 1143) => x"00", (0 + 1144) => x"00", (0 + 1145) => x"00", (0 + 1146) => x"00", (0 + 1147) => x"00", (0 + 1148) => x"00", (0 + 1149) => x"00", (0 + 1150) => x"00", (0 + 1151) => x"00", (0 + 1152) => x"00", (0 + 1153) => x"00", (0 + 1154) => x"00", (0 + 1155) => x"00", (0 + 1156) => x"00", (0 + 1157) => x"00", (0 + 1158) => x"00", (0 + 1159) => x"00", (0 + 1160) => x"00", (0 + 1161) => x"00", (0 + 1162) => x"00", (0 + 1163) => x"00", (0 + 1164) => x"00", (0 + 1165) => x"00", (0 + 1166) => x"00", (0 + 1167) => x"00", (0 + 1168) => x"00", (0 + 1169) => x"00", (0 + 1170) => x"00", (0 + 1171) => x"00", (0 + 1172) => x"00", (0 + 1173) => x"00", (0 + 1174) => x"00", (0 + 1175) => x"00", (0 + 1176) => x"00", (0 + 1177) => x"00", (0 + 1178) => x"00", (0 + 1179) => x"00", (0 + 1180) => x"00", (0 + 1181) => x"00", (0 + 1182) => x"00", (0 + 1183) => x"00", (0 + 1184) => x"00", (0 + 1185) => x"00", (0 + 1186) => x"00", (0 + 1187) => x"00", (0 + 1188) => x"00", (0 + 1189) => x"00", (0 + 1190) => x"00", (0 + 1191) => x"00", (0 + 1192) => x"00", (0 + 1193) => x"00", (0 + 1194) => x"00", (0 + 1195) => x"00", (0 + 1196) => x"00", (0 + 1197) => x"00", (0 + 1198) => x"00", (0 + 1199) => x"00", (0 + 1200) => x"00", (0 + 1201) => x"00", (0 + 1202) => x"00", (0 + 1203) => x"00", (0 + 1204) => x"00", (0 + 1205) => x"00", (0 + 1206) => x"00", (0 + 1207) => x"00", (0 + 1208) => x"00", (0 + 1209) => x"00", (0 + 1210) => x"00", (0 + 1211) => x"00", (0 + 1212) => x"00", (0 + 1213) => x"00", (0 + 1214) => x"00", (0 + 1215) => x"00", (0 + 1216) => x"00", (0 + 1217) => x"00", (0 + 1218) => x"00", (0 + 1219) => x"00", (0 + 1220) => x"00", (0 + 1221) => x"00", (0 + 1222) => x"00", (0 + 1223) => x"00", (0 + 1224) => x"00", (0 + 1225) => x"00", (0 + 1226) => x"00", (0 + 1227) => x"00", (0 + 1228) => x"00", (0 + 1229) => x"00", (0 + 1230) => x"00", (0 + 1231) => x"00", (0 + 1232) => x"00", (0 + 1233) => x"00", (0 + 1234) => x"00", (0 + 1235) => x"00", (0 + 1236) => x"00", (0 + 1237) => x"00", (0 + 1238) => x"00", (0 + 1239) => x"00", (0 + 1240) => x"00", (0 + 1241) => x"00", (0 + 1242) => x"00", (0 + 1243) => x"00", (0 + 1244) => x"00", (0 + 1245) => x"00", (0 + 1246) => x"00", (0 + 1247) => x"00", (0 + 1248) => x"00", (0 + 1249) => x"00", (0 + 1250) => x"00", (0 + 1251) => x"00", (0 + 1252) => x"00", (0 + 1253) => x"00", (0 + 1254) => x"00", (0 + 1255) => x"00", (0 + 1256) => x"00", (0 + 1257) => x"00", (0 + 1258) => x"00", (0 + 1259) => x"00", (0 + 1260) => x"00", (0 + 1261) => x"00", (0 + 1262) => x"00", (0 + 1263) => x"00", (0 + 1264) => x"00", (0 + 1265) => x"00", (0 + 1266) => x"00", (0 + 1267) => x"00", (0 + 1268) => x"00", (0 + 1269) => x"00", (0 + 1270) => x"00", (0 + 1271) => x"00", (0 + 1272) => x"00", (0 + 1273) => x"00", (0 + 1274) => x"00", (0 + 1275) => x"00", (0 + 1276) => x"00", (0 + 1277) => x"00", (0 + 1278) => x"00", (0 + 1279) => x"00", (0 + 1280) => x"00", (0 + 1281) => x"00", (0 + 1282) => x"00", (0 + 1283) => x"00", (0 + 1284) => x"00", (0 + 1285) => x"00", (0 + 1286) => x"00", (0 + 1287) => x"00", (0 + 1288) => x"00", (0 + 1289) => x"00", (0 + 1290) => x"00", (0 + 1291) => x"00", (0 + 1292) => x"00", (0 + 1293) => x"00", (0 + 1294) => x"00", (0 + 1295) => x"00", (0 + 1296) => x"00", (0 + 1297) => x"00", (0 + 1298) => x"00", (0 + 1299) => x"00", (0 + 1300) => x"00", (0 + 1301) => x"00", (0 + 1302) => x"00", (0 + 1303) => x"00", (0 + 1304) => x"00", (0 + 1305) => x"00", (0 + 1306) => x"00", (0 + 1307) => x"00", (0 + 1308) => x"00", (0 + 1309) => x"00", (0 + 1310) => x"00", (0 + 1311) => x"00", (0 + 1312) => x"00", (0 + 1313) => x"00", (0 + 1314) => x"00", (0 + 1315) => x"00", (0 + 1316) => x"00", (0 + 1317) => x"00", (0 + 1318) => x"00", (0 + 1319) => x"00", (0 + 1320) => x"00", (0 + 1321) => x"00", (0 + 1322) => x"00", (0 + 1323) => x"00", (0 + 1324) => x"00", (0 + 1325) => x"00", (0 + 1326) => x"00", (0 + 1327) => x"00", (0 + 1328) => x"00", (0 + 1329) => x"00", (0 + 1330) => x"00", (0 + 1331) => x"00", (0 + 1332) => x"00", (0 + 1333) => x"00", (0 + 1334) => x"00", (0 + 1335) => x"00", (0 + 1336) => x"00", (0 + 1337) => x"00", (0 + 1338) => x"00", (0 + 1339) => x"00", (0 + 1340) => x"00", (0 + 1341) => x"00", (0 + 1342) => x"00", (0 + 1343) => x"00", (0 + 1344) => x"00", (0 + 1345) => x"00", (0 + 1346) => x"00", (0 + 1347) => x"00", (0 + 1348) => x"00", (0 + 1349) => x"00", (0 + 1350) => x"00", (0 + 1351) => x"00", (0 + 1352) => x"00", (0 + 1353) => x"00", (0 + 1354) => x"00", (0 + 1355) => x"00", (0 + 1356) => x"00", (0 + 1357) => x"00", (0 + 1358) => x"00", (0 + 1359) => x"00", (0 + 1360) => x"00", (0 + 1361) => x"00", (0 + 1362) => x"00", (0 + 1363) => x"00", (0 + 1364) => x"00", (0 + 1365) => x"00", (0 + 1366) => x"00", (0 + 1367) => x"00", (0 + 1368) => x"00", (0 + 1369) => x"00", (0 + 1370) => x"00", (0 + 1371) => x"00", (0 + 1372) => x"00", (0 + 1373) => x"00", (0 + 1374) => x"00", (0 + 1375) => x"00", (0 + 1376) => x"00", (0 + 1377) => x"00", (0 + 1378) => x"00", (0 + 1379) => x"00", (0 + 1380) => x"00", (0 + 1381) => x"00", (0 + 1382) => x"00", (0 + 1383) => x"00", (0 + 1384) => x"00", (0 + 1385) => x"00", (0 + 1386) => x"00", (0 + 1387) => x"00", (0 + 1388) => x"00", (0 + 1389) => x"00", (0 + 1390) => x"00", (0 + 1391) => x"00", (0 + 1392) => x"00", (0 + 1393) => x"00", (0 + 1394) => x"00", (0 + 1395) => x"00", (0 + 1396) => x"00", (0 + 1397) => x"00", (0 + 1398) => x"00", (0 + 1399) => x"00", (0 + 1400) => x"00", (0 + 1401) => x"00", (0 + 1402) => x"00", (0 + 1403) => x"00", (0 + 1404) => x"00", (0 + 1405) => x"00", (0 + 1406) => x"00", (0 + 1407) => x"00", (0 + 1408) => x"00", (0 + 1409) => x"00", (0 + 1410) => x"00", (0 + 1411) => x"00", (0 + 1412) => x"00", (0 + 1413) => x"00", (0 + 1414) => x"00", (0 + 1415) => x"00", (0 + 1416) => x"00", (0 + 1417) => x"00", (0 + 1418) => x"00", (0 + 1419) => x"00", (0 + 1420) => x"00", (0 + 1421) => x"00", (0 + 1422) => x"00", (0 + 1423) => x"00", (0 + 1424) => x"00", (0 + 1425) => x"00", (0 + 1426) => x"00", (0 + 1427) => x"00", (0 + 1428) => x"00", (0 + 1429) => x"00", (0 + 1430) => x"00", (0 + 1431) => x"00", (0 + 1432) => x"00", (0 + 1433) => x"00", (0 + 1434) => x"00", (0 + 1435) => x"00", (0 + 1436) => x"00", (0 + 1437) => x"00", (0 + 1438) => x"00", (0 + 1439) => x"00", (0 + 1440) => x"00", (0 + 1441) => x"00", (0 + 1442) => x"00", (0 + 1443) => x"00", (0 + 1444) => x"00", (0 + 1445) => x"00", (0 + 1446) => x"00", (0 + 1447) => x"00", (0 + 1448) => x"00", (0 + 1449) => x"00", (0 + 1450) => x"00", (0 + 1451) => x"00", (0 + 1452) => x"00", (0 + 1453) => x"00", (0 + 1454) => x"00", (0 + 1455) => x"00", (0 + 1456) => x"00", (0 + 1457) => x"00", (0 + 1458) => x"00", (0 + 1459) => x"00", (0 + 1460) => x"00", (0 + 1461) => x"00", (0 + 1462) => x"00", (0 + 1463) => x"00", (0 + 1464) => x"00", (0 + 1465) => x"00", (0 + 1466) => x"00", (0 + 1467) => x"00", (0 + 1468) => x"00", (0 + 1469) => x"00", (0 + 1470) => x"00", (0 + 1471) => x"00", (0 + 1472) => x"00", (0 + 1473) => x"00", (0 + 1474) => x"00", (0 + 1475) => x"00", (0 + 1476) => x"00", (0 + 1477) => x"00", (0 + 1478) => x"00", (0 + 1479) => x"00", (0 + 1480) => x"00", (0 + 1481) => x"00", (0 + 1482) => x"00", (0 + 1483) => x"00", (0 + 1484) => x"00", (0 + 1485) => x"00", (0 + 1486) => x"00", (0 + 1487) => x"00", (0 + 1488) => x"00", (0 + 1489) => x"00", (0 + 1490) => x"00", (0 + 1491) => x"00", (0 + 1492) => x"00", (0 + 1493) => x"00", (0 + 1494) => x"00", (0 + 1495) => x"00", (0 + 1496) => x"00", (0 + 1497) => x"00", (0 + 1498) => x"00", (0 + 1499) => x"00", (0 + 1500) => x"00", (0 + 1501) => x"00", (0 + 1502) => x"00", (0 + 1503) => x"00", (0 + 1504) => x"00", (0 + 1505) => x"00", (0 + 1506) => x"00", (0 + 1507) => x"00", (0 + 1508) => x"00", (0 + 1509) => x"00", (0 + 1510) => x"00", (0 + 1511) => x"00", (0 + 1512) => x"00", (0 + 1513) => x"00", (0 + 1514) => x"00", (0 + 1515) => x"00", (0 + 1516) => x"00", (0 + 1517) => x"00", (0 + 1518) => x"00", (0 + 1519) => x"00", (0 + 1520) => x"00", (0 + 1521) => x"00", (0 + 1522) => x"00", (0 + 1523) => x"00", (0 + 1524) => x"00", (0 + 1525) => x"00", (0 + 1526) => x"00", (0 + 1527) => x"00", (0 + 1528) => x"00", (0 + 1529) => x"00", (0 + 1530) => x"00", (0 + 1531) => x"00", (0 + 1532) => x"00", (0 + 1533) => x"00", (0 + 1534) => x"00", (0 + 1535) => x"00", (0 + 1536) => x"00", (0 + 1537) => x"00", (0 + 1538) => x"00", (0 + 1539) => x"00", (0 + 1540) => x"00", (0 + 1541) => x"00", (0 + 1542) => x"00", (0 + 1543) => x"00", (0 + 1544) => x"00", (0 + 1545) => x"00", (0 + 1546) => x"00", (0 + 1547) => x"00", (0 + 1548) => x"00", (0 + 1549) => x"00", (0 + 1550) => x"00", (0 + 1551) => x"00", (0 + 1552) => x"00", (0 + 1553) => x"00", (0 + 1554) => x"00", (0 + 1555) => x"00", (0 + 1556) => x"00", (0 + 1557) => x"00", (0 + 1558) => x"00", (0 + 1559) => x"00", (0 + 1560) => x"00", (0 + 1561) => x"00", (0 + 1562) => x"00", (0 + 1563) => x"00", (0 + 1564) => x"00", (0 + 1565) => x"00", (0 + 1566) => x"00", (0 + 1567) => x"00", (0 + 1568) => x"00", (0 + 1569) => x"00", (0 + 1570) => x"00", (0 + 1571) => x"00", (0 + 1572) => x"00", (0 + 1573) => x"00", (0 + 1574) => x"00", (0 + 1575) => x"00", (0 + 1576) => x"00", (0 + 1577) => x"00", (0 + 1578) => x"00", (0 + 1579) => x"00", (0 + 1580) => x"00", (0 + 1581) => x"00", (0 + 1582) => x"00", (0 + 1583) => x"00", (0 + 1584) => x"00", (0 + 1585) => x"00", (0 + 1586) => x"00", (0 + 1587) => x"00", (0 + 1588) => x"00", (0 + 1589) => x"00", (0 + 1590) => x"00", (0 + 1591) => x"00", (0 + 1592) => x"00", (0 + 1593) => x"00", (0 + 1594) => x"00", (0 + 1595) => x"00", (0 + 1596) => x"00", (0 + 1597) => x"00", (0 + 1598) => x"00", (0 + 1599) => x"00", (0 + 1600) => x"00", (0 + 1601) => x"00", (0 + 1602) => x"00", (0 + 1603) => x"00", (0 + 1604) => x"00", (0 + 1605) => x"00", (0 + 1606) => x"00", (0 + 1607) => x"00", (0 + 1608) => x"00", (0 + 1609) => x"00", (0 + 1610) => x"00", (0 + 1611) => x"00", (0 + 1612) => x"00", (0 + 1613) => x"00", (0 + 1614) => x"00", (0 + 1615) => x"00", (0 + 1616) => x"00", (0 + 1617) => x"00", (0 + 1618) => x"00", (0 + 1619) => x"00", (0 + 1620) => x"00", (0 + 1621) => x"00", (0 + 1622) => x"00", (0 + 1623) => x"00", (0 + 1624) => x"00", (0 + 1625) => x"00", (0 + 1626) => x"00", (0 + 1627) => x"00", (0 + 1628) => x"00", (0 + 1629) => x"00", (0 + 1630) => x"00", (0 + 1631) => x"00", (0 + 1632) => x"00", (0 + 1633) => x"00", (0 + 1634) => x"00", (0 + 1635) => x"00", (0 + 1636) => x"00", (0 + 1637) => x"00", (0 + 1638) => x"00", (0 + 1639) => x"00", (0 + 1640) => x"00", (0 + 1641) => x"00", (0 + 1642) => x"00", (0 + 1643) => x"00", (0 + 1644) => x"00", (0 + 1645) => x"00", (0 + 1646) => x"00", (0 + 1647) => x"00", (0 + 1648) => x"00", (0 + 1649) => x"00", (0 + 1650) => x"00", (0 + 1651) => x"00", (0 + 1652) => x"00", (0 + 1653) => x"00", (0 + 1654) => x"00", (0 + 1655) => x"00", (0 + 1656) => x"00", (0 + 1657) => x"00", (0 + 1658) => x"00", (0 + 1659) => x"00", (0 + 1660) => x"00", (0 + 1661) => x"00", (0 + 1662) => x"00", (0 + 1663) => x"00", (0 + 1664) => x"00", (0 + 1665) => x"00", (0 + 1666) => x"00", (0 + 1667) => x"00", (0 + 1668) => x"00", (0 + 1669) => x"00", (0 + 1670) => x"00", (0 + 1671) => x"00", (0 + 1672) => x"00", (0 + 1673) => x"00", (0 + 1674) => x"00", (0 + 1675) => x"00", (0 + 1676) => x"00", (0 + 1677) => x"00", (0 + 1678) => x"00", (0 + 1679) => x"00", (0 + 1680) => x"00", (0 + 1681) => x"00", (0 + 1682) => x"00", (0 + 1683) => x"00", (0 + 1684) => x"00", (0 + 1685) => x"00", (0 + 1686) => x"00", (0 + 1687) => x"00", (0 + 1688) => x"00", (0 + 1689) => x"00", (0 + 1690) => x"00", (0 + 1691) => x"00", (0 + 1692) => x"00", (0 + 1693) => x"00", (0 + 1694) => x"00", (0 + 1695) => x"00", (0 + 1696) => x"00", (0 + 1697) => x"00", (0 + 1698) => x"00", (0 + 1699) => x"00", (0 + 1700) => x"00", (0 + 1701) => x"00", (0 + 1702) => x"00", (0 + 1703) => x"00", (0 + 1704) => x"00", (0 + 1705) => x"00", (0 + 1706) => x"00", (0 + 1707) => x"00", (0 + 1708) => x"00", (0 + 1709) => x"00", (0 + 1710) => x"00", (0 + 1711) => x"00", (0 + 1712) => x"00", (0 + 1713) => x"00", (0 + 1714) => x"00", (0 + 1715) => x"00", (0 + 1716) => x"00", (0 + 1717) => x"00", (0 + 1718) => x"00", (0 + 1719) => x"00", (0 + 1720) => x"00", (0 + 1721) => x"00", (0 + 1722) => x"00", (0 + 1723) => x"00", (0 + 1724) => x"00", (0 + 1725) => x"00", (0 + 1726) => x"00", (0 + 1727) => x"00", (0 + 1728) => x"00", (0 + 1729) => x"00", (0 + 1730) => x"00", (0 + 1731) => x"00", (0 + 1732) => x"00", (0 + 1733) => x"00", (0 + 1734) => x"00", (0 + 1735) => x"00", (0 + 1736) => x"00", (0 + 1737) => x"00", (0 + 1738) => x"00", (0 + 1739) => x"00", (0 + 1740) => x"00", (0 + 1741) => x"00", (0 + 1742) => x"00", (0 + 1743) => x"00", (0 + 1744) => x"00", (0 + 1745) => x"00", (0 + 1746) => x"00", (0 + 1747) => x"00", (0 + 1748) => x"00", (0 + 1749) => x"00", (0 + 1750) => x"00", (0 + 1751) => x"00", (0 + 1752) => x"00", (0 + 1753) => x"00", (0 + 1754) => x"00", (0 + 1755) => x"00", (0 + 1756) => x"00", (0 + 1757) => x"00", (0 + 1758) => x"00", (0 + 1759) => x"00", (0 + 1760) => x"00", (0 + 1761) => x"00", (0 + 1762) => x"00", (0 + 1763) => x"00", (0 + 1764) => x"00", (0 + 1765) => x"00", (0 + 1766) => x"00", (0 + 1767) => x"00", (0 + 1768) => x"00", (0 + 1769) => x"00", (0 + 1770) => x"00", (0 + 1771) => x"00", (0 + 1772) => x"00", (0 + 1773) => x"00", (0 + 1774) => x"00", (0 + 1775) => x"00", (0 + 1776) => x"00", (0 + 1777) => x"00", (0 + 1778) => x"00", (0 + 1779) => x"00", (0 + 1780) => x"00", (0 + 1781) => x"00", (0 + 1782) => x"00", (0 + 1783) => x"00", (0 + 1784) => x"00", (0 + 1785) => x"00", (0 + 1786) => x"00", (0 + 1787) => x"00", (0 + 1788) => x"00", (0 + 1789) => x"00", (0 + 1790) => x"00", (0 + 1791) => x"00", (0 + 1792) => x"00", (0 + 1793) => x"00", (0 + 1794) => x"00", (0 + 1795) => x"00", (0 + 1796) => x"00", (0 + 1797) => x"00", (0 + 1798) => x"00", (0 + 1799) => x"00", (0 + 1800) => x"00", (0 + 1801) => x"00", (0 + 1802) => x"00", (0 + 1803) => x"00", (0 + 1804) => x"00", (0 + 1805) => x"00", (0 + 1806) => x"00", (0 + 1807) => x"00", (0 + 1808) => x"00", (0 + 1809) => x"00", (0 + 1810) => x"00", (0 + 1811) => x"00", (0 + 1812) => x"00", (0 + 1813) => x"00", (0 + 1814) => x"00", (0 + 1815) => x"00", (0 + 1816) => x"00", (0 + 1817) => x"00", (0 + 1818) => x"00", (0 + 1819) => x"00", (0 + 1820) => x"00", (0 + 1821) => x"00", (0 + 1822) => x"00", (0 + 1823) => x"00", (0 + 1824) => x"00", (0 + 1825) => x"00", (0 + 1826) => x"00", (0 + 1827) => x"00", (0 + 1828) => x"00", (0 + 1829) => x"00", (0 + 1830) => x"00", (0 + 1831) => x"00", (0 + 1832) => x"00", (0 + 1833) => x"00", (0 + 1834) => x"00", (0 + 1835) => x"00", (0 + 1836) => x"00", (0 + 1837) => x"00", (0 + 1838) => x"00", (0 + 1839) => x"00", (0 + 1840) => x"00", (0 + 1841) => x"00", (0 + 1842) => x"00", (0 + 1843) => x"00", (0 + 1844) => x"00", (0 + 1845) => x"00", (0 + 1846) => x"00", (0 + 1847) => x"00", (0 + 1848) => x"00", (0 + 1849) => x"00", (0 + 1850) => x"00", (0 + 1851) => x"00", (0 + 1852) => x"00", (0 + 1853) => x"00", (0 + 1854) => x"00", (0 + 1855) => x"00", (0 + 1856) => x"00", (0 + 1857) => x"00", (0 + 1858) => x"00", (0 + 1859) => x"00", (0 + 1860) => x"00", (0 + 1861) => x"00", (0 + 1862) => x"00", (0 + 1863) => x"00", (0 + 1864) => x"00", (0 + 1865) => x"00", (0 + 1866) => x"00", (0 + 1867) => x"00", (0 + 1868) => x"00", (0 + 1869) => x"00", (0 + 1870) => x"00", (0 + 1871) => x"00", (0 + 1872) => x"00", (0 + 1873) => x"00", (0 + 1874) => x"00", (0 + 1875) => x"00", (0 + 1876) => x"00", (0 + 1877) => x"00", (0 + 1878) => x"00", (0 + 1879) => x"00", (0 + 1880) => x"00", (0 + 1881) => x"00", (0 + 1882) => x"00", (0 + 1883) => x"00", (0 + 1884) => x"00", (0 + 1885) => x"00", (0 + 1886) => x"00", (0 + 1887) => x"00", (0 + 1888) => x"00", (0 + 1889) => x"00", (0 + 1890) => x"00", (0 + 1891) => x"00", (0 + 1892) => x"00", (0 + 1893) => x"00", (0 + 1894) => x"00", (0 + 1895) => x"00", (0 + 1896) => x"00", (0 + 1897) => x"00", (0 + 1898) => x"00", (0 + 1899) => x"00", (0 + 1900) => x"00", (0 + 1901) => x"00", (0 + 1902) => x"00", (0 + 1903) => x"00", (0 + 1904) => x"00", (0 + 1905) => x"00", (0 + 1906) => x"00", (0 + 1907) => x"00", (0 + 1908) => x"00", (0 + 1909) => x"00", (0 + 1910) => x"00", (0 + 1911) => x"00", (0 + 1912) => x"00", (0 + 1913) => x"00", (0 + 1914) => x"00", (0 + 1915) => x"00", (0 + 1916) => x"00", (0 + 1917) => x"00", (0 + 1918) => x"00", (0 + 1919) => x"00", (0 + 1920) => x"00", (0 + 1921) => x"00", (0 + 1922) => x"00", (0 + 1923) => x"00", (0 + 1924) => x"00", (0 + 1925) => x"00", (0 + 1926) => x"00", (0 + 1927) => x"00", (0 + 1928) => x"00", (0 + 1929) => x"00", (0 + 1930) => x"00", (0 + 1931) => x"00", (0 + 1932) => x"00", (0 + 1933) => x"00", (0 + 1934) => x"00", (0 + 1935) => x"00", (0 + 1936) => x"00", (0 + 1937) => x"00", (0 + 1938) => x"00", (0 + 1939) => x"00", (0 + 1940) => x"00", (0 + 1941) => x"00", (0 + 1942) => x"00", (0 + 1943) => x"00", (0 + 1944) => x"00", (0 + 1945) => x"00", (0 + 1946) => x"00", (0 + 1947) => x"00", (0 + 1948) => x"00", (0 + 1949) => x"00", (0 + 1950) => x"00", (0 + 1951) => x"00", (0 + 1952) => x"00", (0 + 1953) => x"00", (0 + 1954) => x"00", (0 + 1955) => x"00", (0 + 1956) => x"00", (0 + 1957) => x"00", (0 + 1958) => x"00", (0 + 1959) => x"00", (0 + 1960) => x"00", (0 + 1961) => x"00", (0 + 1962) => x"00", (0 + 1963) => x"00", (0 + 1964) => x"00", (0 + 1965) => x"00", (0 + 1966) => x"00", (0 + 1967) => x"00", (0 + 1968) => x"00", (0 + 1969) => x"00", (0 + 1970) => x"00", (0 + 1971) => x"00", (0 + 1972) => x"00", (0 + 1973) => x"00", (0 + 1974) => x"00", (0 + 1975) => x"00", (0 + 1976) => x"00", (0 + 1977) => x"00", (0 + 1978) => x"00", (0 + 1979) => x"00", (0 + 1980) => x"00", (0 + 1981) => x"00", (0 + 1982) => x"00", (0 + 1983) => x"00", (0 + 1984) => x"00", (0 + 1985) => x"00", (0 + 1986) => x"00", (0 + 1987) => x"00", (0 + 1988) => x"00", (0 + 1989) => x"00", (0 + 1990) => x"00", (0 + 1991) => x"00", (0 + 1992) => x"00", (0 + 1993) => x"00", (0 + 1994) => x"00", (0 + 1995) => x"00", (0 + 1996) => x"00", (0 + 1997) => x"00", (0 + 1998) => x"00", (0 + 1999) => x"00", (0 + 2000) => x"00", (0 + 2001) => x"00", (0 + 2002) => x"00", (0 + 2003) => x"00", (0 + 2004) => x"00", (0 + 2005) => x"00", (0 + 2006) => x"00", (0 + 2007) => x"00", (0 + 2008) => x"00", (0 + 2009) => x"00", (0 + 2010) => x"00", (0 + 2011) => x"00", (0 + 2012) => x"00", (0 + 2013) => x"00", (0 + 2014) => x"00", (0 + 2015) => x"00", (0 + 2016) => x"00", (0 + 2017) => x"00", (0 + 2018) => x"00", (0 + 2019) => x"00", (0 + 2020) => x"00", (0 + 2021) => x"00", (0 + 2022) => x"00", (0 + 2023) => x"00", (0 + 2024) => x"00", (0 + 2025) => x"00", (0 + 2026) => x"00", (0 + 2027) => x"00", (0 + 2028) => x"00", (0 + 2029) => x"00", (0 + 2030) => x"00", (0 + 2031) => x"00", (0 + 2032) => x"00", (0 + 2033) => x"00", (0 + 2034) => x"00", (0 + 2035) => x"00", (0 + 2036) => x"00", (0 + 2037) => x"00", (0 + 2038) => x"00", (0 + 2039) => x"00", (0 + 2040) => x"00", (0 + 2041) => x"00", (0 + 2042) => x"00", (0 + 2043) => x"00", (0 + 2044) => x"00", (0 + 2045) => x"00", (0 + 2046) => x"00", (0 + 2047) => x"00", 
                                others => ( others => '0')
                            );
    
    signal read_address : std_logic_vector( 11 downto 0 );
begin

    process ( clock )
    begin
        if ( rising_edge( clock ) ) then
            if( we = '1' ) then
                sys_RAM( to_integer( unsigned( address ))) <= dataIn;
            end if;
            
            read_address <= address;
        end if;
    end process;

    dataOut <= sys_RAM( to_integer( unsigned( read_address )));
end Behavioral;
